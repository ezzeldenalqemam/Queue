<svg width="116" height="33" viewBox="0 0 116 33" fill="none" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink">
<rect width="32" height="32" transform="translate(0.664062 0.980469)" fill="url(#pattern0_1_3640)"/>
<path d="M47.8041 21.9205C48.0841 22.3031 48.3734 22.6065 48.6721 22.8305C48.9707 23.0545 49.2834 23.1665 49.6101 23.1665C49.8621 23.1665 50.1421 23.0918 50.4501 22.9425C50.7581 22.8025 51.0661 22.6065 51.3741 22.3545L52.1021 23.5725C51.7287 23.9178 51.2994 24.1838 50.8141 24.3705C50.3287 24.5665 49.8527 24.6645 49.3861 24.6645C48.7421 24.6645 48.1447 24.4685 47.5941 24.0765C47.0434 23.6938 46.5861 23.1618 46.2221 22.4805L47.8041 21.9205ZM46.3201 12.5685C47.0574 12.5685 47.7434 12.6945 48.3781 12.9465C49.0127 13.1985 49.5634 13.5531 50.0301 14.0105C50.5061 14.4678 50.8747 14.9998 51.1361 15.6065C51.4067 16.2038 51.5421 16.8571 51.5421 17.5665C51.5421 18.2665 51.4067 18.9245 51.1361 19.5405C50.8747 20.1565 50.5061 20.6931 50.0301 21.1505C49.5634 21.6078 49.0127 21.9671 48.3781 22.2285C47.7434 22.4805 47.0574 22.6065 46.3201 22.6065C45.5827 22.6065 44.8967 22.4805 44.2621 22.2285C43.6367 21.9671 43.0861 21.6078 42.6101 21.1505C42.1341 20.6931 41.7607 20.1611 41.4901 19.5545C41.2287 18.9385 41.0981 18.2758 41.0981 17.5665C41.0981 16.8571 41.2287 16.1991 41.4901 15.5925C41.7607 14.9858 42.1341 14.4585 42.6101 14.0105C43.0861 13.5531 43.6367 13.1985 44.2621 12.9465C44.8967 12.6945 45.5827 12.5685 46.3201 12.5685ZM46.3481 14.1505C45.8907 14.1505 45.4614 14.2391 45.0601 14.4165C44.6587 14.5845 44.3041 14.8271 43.9961 15.1445C43.6881 15.4525 43.4454 15.8118 43.2681 16.2225C43.1001 16.6331 43.0161 17.0811 43.0161 17.5665C43.0161 18.0518 43.1047 18.5045 43.2821 18.9245C43.4594 19.3351 43.7021 19.6991 44.0101 20.0165C44.3181 20.3338 44.6727 20.5811 45.0741 20.7585C45.4754 20.9358 45.9001 21.0245 46.3481 21.0245C46.7961 21.0245 47.2161 20.9358 47.6081 20.7585C48.0094 20.5811 48.3594 20.3338 48.6581 20.0165C48.9567 19.6991 49.1901 19.3351 49.3581 18.9245C49.5354 18.5045 49.6241 18.0518 49.6241 17.5665C49.6241 17.0811 49.5354 16.6331 49.3581 16.2225C49.1901 15.8118 48.9567 15.4525 48.6581 15.1445C48.3594 14.8271 48.0094 14.5845 47.6081 14.4165C47.2161 14.2391 46.7961 14.1505 46.3481 14.1505ZM54.8238 19.1765C54.8238 19.7178 54.9638 20.1471 55.2438 20.4645C55.5331 20.7725 55.9298 20.9265 56.4338 20.9265C57.0218 20.9078 57.4791 20.6885 57.8058 20.2685C58.1418 19.8485 58.3098 19.3211 58.3098 18.6865H58.7858C58.7858 19.5918 58.6598 20.3291 58.4078 20.8985C58.1558 21.4585 57.8011 21.8738 57.3438 22.1445C56.8864 22.4058 56.3404 22.5411 55.7058 22.5505C55.1458 22.5505 54.6604 22.4338 54.2498 22.2005C53.8484 21.9671 53.5358 21.6358 53.3118 21.2065C53.0971 20.7678 52.9898 20.2545 52.9898 19.6665V15.0185H54.8238V19.1765ZM58.3098 15.0185H60.1438V22.4805H58.3098V15.0185ZM67.4693 18.1825C67.4506 17.7905 67.3619 17.4591 67.2033 17.1885C67.0446 16.9085 66.8206 16.6938 66.5313 16.5445C66.2513 16.3858 65.9293 16.3065 65.5653 16.3065C65.1453 16.3065 64.7813 16.4045 64.4733 16.6005C64.1653 16.7965 63.9226 17.0718 63.7453 17.4265C63.5773 17.7811 63.4933 18.1918 63.4933 18.6585C63.4933 19.1718 63.5866 19.6151 63.7733 19.9885C63.9693 20.3618 64.2353 20.6511 64.5713 20.8565C64.9073 21.0525 65.2946 21.1505 65.7333 21.1505C66.5266 21.1505 67.2033 20.8658 67.7633 20.2965L68.7293 21.2625C68.3559 21.6731 67.9033 21.9905 67.3713 22.2145C66.8393 22.4385 66.2466 22.5505 65.5933 22.5505C64.8093 22.5505 64.1279 22.3918 63.5493 22.0745C62.9799 21.7478 62.5319 21.3045 62.2052 20.7445C61.8879 20.1751 61.7293 19.5125 61.7293 18.7565C61.7293 18.0005 61.8879 17.3378 62.2052 16.7685C62.5319 16.1991 62.9799 15.7558 63.5493 15.4385C64.1279 15.1211 64.7906 14.9578 65.5373 14.9485C66.4239 14.9485 67.1379 15.1305 67.6793 15.4945C68.2299 15.8585 68.6219 16.3718 68.8553 17.0345C69.0886 17.6878 69.1726 18.4671 69.1073 19.3725H63.2273V18.1825H67.4693ZM72.2964 19.1765C72.2964 19.7178 72.4364 20.1471 72.7164 20.4645C73.0057 20.7725 73.4024 20.9265 73.9064 20.9265C74.4944 20.9078 74.9517 20.6885 75.2784 20.2685C75.6144 19.8485 75.7824 19.3211 75.7824 18.6865H76.2584C76.2584 19.5918 76.1324 20.3291 75.8804 20.8985C75.6284 21.4585 75.2737 21.8738 74.8164 22.1445C74.3591 22.4058 73.8131 22.5411 73.1784 22.5505C72.6184 22.5505 72.1331 22.4338 71.7224 22.2005C71.3211 21.9671 71.0084 21.6358 70.7844 21.2065C70.5697 20.7678 70.4624 20.2545 70.4624 19.6665V15.0185H72.2964V19.1765ZM75.7824 15.0185H77.6164V22.4805H75.7824V15.0185ZM84.9419 18.1825C84.9232 17.7905 84.8346 17.4591 84.6759 17.1885C84.5172 16.9085 84.2932 16.6938 84.0039 16.5445C83.7239 16.3858 83.4019 16.3065 83.0379 16.3065C82.6179 16.3065 82.2539 16.4045 81.9459 16.6005C81.6379 16.7965 81.3952 17.0718 81.2179 17.4265C81.0499 17.7811 80.9659 18.1918 80.9659 18.6585C80.9659 19.1718 81.0592 19.6151 81.2459 19.9885C81.4419 20.3618 81.7079 20.6511 82.0439 20.8565C82.3799 21.0525 82.7672 21.1505 83.2059 21.1505C83.9992 21.1505 84.6759 20.8658 85.2359 20.2965L86.2019 21.2625C85.8286 21.6731 85.3759 21.9905 84.8439 22.2145C84.3119 22.4385 83.7192 22.5505 83.0659 22.5505C82.2819 22.5505 81.6006 22.3918 81.0219 22.0745C80.4526 21.7478 80.0046 21.3045 79.6779 20.7445C79.3606 20.1751 79.2019 19.5125 79.2019 18.7565C79.2019 18.0005 79.3606 17.3378 79.6779 16.7685C80.0046 16.1991 80.4526 15.7558 81.0219 15.4385C81.6006 15.1211 82.2632 14.9578 83.0099 14.9485C83.8966 14.9485 84.6106 15.1305 85.1519 15.4945C85.7026 15.8585 86.0946 16.3718 86.3279 17.0345C86.5612 17.6878 86.6452 18.4671 86.5799 19.3725H80.6999V18.1825H84.9419ZM96.3565 14.9485C97.0658 14.9485 97.6865 15.1071 98.2185 15.4245C98.7505 15.7418 99.1612 16.1898 99.4505 16.7685C99.7492 17.3378 99.8985 18.0051 99.8985 18.7705C99.8985 19.5171 99.7538 20.1751 99.4645 20.7445C99.1752 21.3045 98.7645 21.7478 98.2325 22.0745C97.7098 22.3918 97.0938 22.5505 96.3845 22.5505C95.7218 22.5505 95.1525 22.4011 94.6765 22.1025C94.2005 21.7945 93.8365 21.3558 93.5845 20.7865C93.3325 20.2171 93.2065 19.5451 93.2065 18.7705C93.2065 17.9678 93.3278 17.2818 93.5705 16.7125C93.8225 16.1431 94.1865 15.7091 94.6625 15.4105C95.1385 15.1025 95.7032 14.9485 96.3565 14.9485ZM95.9505 16.3905C95.5398 16.3905 95.1712 16.4931 94.8445 16.6985C94.5272 16.8945 94.2798 17.1698 94.1025 17.5245C93.9252 17.8698 93.8365 18.2711 93.8365 18.7285C93.8365 19.1858 93.9252 19.5918 94.1025 19.9465C94.2798 20.3011 94.5272 20.5765 94.8445 20.7725C95.1712 20.9685 95.5398 21.0665 95.9505 21.0665C96.3705 21.0665 96.7345 20.9685 97.0425 20.7725C97.3598 20.5671 97.6072 20.2918 97.7845 19.9465C97.9618 19.5918 98.0505 19.1858 98.0505 18.7285C98.0505 18.2711 97.9618 17.8698 97.7845 17.5245C97.6072 17.1698 97.3598 16.8945 97.0425 16.6985C96.7345 16.4931 96.3705 16.3905 95.9505 16.3905ZM92.0165 12.0925H93.8365V22.4805H92.0165V12.0925ZM104.752 14.9485C105.526 14.9485 106.208 15.1071 106.796 15.4245C107.393 15.7418 107.855 16.1851 108.182 16.7545C108.518 17.3238 108.686 17.9865 108.686 18.7425C108.686 19.4985 108.518 20.1611 108.182 20.7305C107.855 21.2998 107.393 21.7478 106.796 22.0745C106.208 22.3918 105.526 22.5505 104.752 22.5505C103.968 22.5505 103.277 22.3918 102.68 22.0745C102.082 21.7478 101.616 21.2998 101.28 20.7305C100.953 20.1611 100.79 19.4985 100.79 18.7425C100.79 17.9865 100.953 17.3238 101.28 16.7545C101.616 16.1851 102.082 15.7418 102.68 15.4245C103.277 15.1071 103.968 14.9485 104.752 14.9485ZM104.752 16.4185C104.332 16.4185 103.958 16.5211 103.632 16.7265C103.314 16.9225 103.067 17.1978 102.89 17.5525C102.712 17.8978 102.624 18.2991 102.624 18.7565C102.624 19.2231 102.712 19.6338 102.89 19.9885C103.067 20.3431 103.314 20.6185 103.632 20.8145C103.958 21.0105 104.332 21.1085 104.752 21.1085C105.162 21.1085 105.526 21.0105 105.844 20.8145C106.161 20.6185 106.408 20.3431 106.586 19.9885C106.763 19.6338 106.852 19.2231 106.852 18.7565C106.852 18.2991 106.763 17.8978 106.586 17.5525C106.408 17.1978 106.161 16.9225 105.844 16.7265C105.526 16.5211 105.162 16.4185 104.752 16.4185ZM112.381 20.0445C112.381 20.4178 112.451 20.6745 112.591 20.8145C112.731 20.9545 112.922 21.0245 113.165 21.0245C113.314 21.0245 113.477 21.0011 113.655 20.9545C113.832 20.8985 114.023 20.8145 114.229 20.7025L114.649 22.0185C114.369 22.1865 114.065 22.3218 113.739 22.4245C113.421 22.5178 113.099 22.5645 112.773 22.5645C112.371 22.5645 112.003 22.4898 111.667 22.3405C111.331 22.1818 111.065 21.9391 110.869 21.6125C110.673 21.2765 110.575 20.8565 110.575 20.3525V13.2545H112.381V20.0445ZM109.525 15.2985H114.523V16.5725H109.525V15.2985Z" fill="white"/>
<defs>
<pattern id="pattern0_1_3640" patternContentUnits="objectBoundingBox" width="1" height="1">
<use xlink:href="#image0_1_3640" transform="translate(0.0786498 0.15625) scale(0.000664741)"/>
</pattern>
<image id="image0_1_3640" width="3365" height="1014" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAADSUAAAP2CAYAAACrSBkYAAAACXBIWXMAAC4jAAAuIwF4pT92AAAgAElEQVR4nOzd/XEbZ5bo4SPV/g/cCAhHQGwEhCMgHQGhCExHICoCUxEIjGCoCAaMwEAEl8wAiAC3eubwDobmF4AG0N3v81Sx7PV6t9DnlcWmqn99Pq1WqwAAeMEgv/bpIb8AAAAAAAAAAAAAgBb5H4cFAK02evbhhxHRf/bPnv87T85acuHziFi88M9nL/zz6Qf+HQAAAAAAAAAAAABgRzYlAUAz9DMoimcbitb/eeTf95zZ1u7X/g/XtzS99vcAAAAAAAAAAAAAwAtESQCwX0+bi9bjovV/dmr+jba+pelpC9N6tPR8MxMAAAAAAAAAAAAAFEGUBADbGzz7Wg+Pzsy1KE/x0sOzr+qfzUofDgAAAAAAAAAAAADdI0oCgNc9RUbP46Pq68Tc2MAy46SnSOl5vAQAAAAAAAAAAAAArSJKAqB0T+HRMP9+lH89LX0wHNTTpqXpC+ESAAAAAAAAAAAAADSOKAmAUjxtPFoPkM6cPi0wzzhpPVSaOjgAAAAAAAAAAAAAjkmUBEDXPI+PBrYe0VGPa4GSWAkAAAAAAAAAAACAgxIlAdBWg/waiY/gvzzmVqX1rwcjAgAAAAAAAAAAAKBOoiQA2mD4wlfPycFG7uM/gdLMViUAAAAAAAAAAAAAdiFKAqBpngdIZ04I9mb+bKOSUAkAAAAAAAAAAACADxElAXBMAiRonvmzSGnmjAAAAAAAAAAAAAB4TpQEwKH0I2KU8dHTX3umD61w/yxSenBsAAAAAAAAAAAAAGUTJQGwL8NnEdKJSUNnPD6LlKaOFgAAAAAAAAAAAKAsoiQA6jJa+7IFCcpz/yxSWvg1AAAAAAAAAAAAANBdoiQAttF/FiCdmSLwzDzjpKlICQAAAAAAAAAAAKB7REkAfET/2SakU1MDNiRSAgAAAAAAAAAAAOgQURIAr6niowsRErAnIiUAAAAAAAAAAACAFhMlAfBkuBYhnZkKcGBPkdJd/hUAAAAAAAAAAACABhMlAZRr8GwbUs+vBaBBfq5tUZo5GAAAAAAAAAAAAIBmESUBlOViLUQ6cfZASzw+26K0cHAAAAAAAAAAAAAAxyVKAui2wVqIdO6sgY6YZ6B0Z4sSAAAAAAAAAAAAwHGIkgC6xzYkoCS2KAEAAAAAAAAAAAAcgSgJoP36GSA9xUg9ZwoU7OdapPTgFwIAAAAAAAAAAADAfoiSANppsBYinTlDgBfNM06qvmZGBAAAAAAAAAAAAFAfURJAewwjYpzbkE6dG8BGHtcCpanRAQAAAAAAAAAAAOxGlATQbE8hUrUR6cRZAdRiuRYo3RkpAAAAAAAAAAAAwOZESQDNc5HbkIRIAPsnUAIAAAAAAAAAAADYgigJoBku1r56zgTgKARKAAAAAAAAAAAAAB8kSgI4nmFEjG1EAmgkgRIAAAAAAAAAAADAG0RJAIclRAJon6dAaRIRU+cHAAAAAAAAAAAAIEoCOIRBhkhjIRJA6z2uBUozxwkAAAAAAAAAAACUSpQEsB/9tRDp1IwBOqkKlG4yUnpwxAAAAAAAAAAAAEBJREkA9aoipIuIODdXgKLc5/akKlBaOHoAAAAAAAAAAACg60RJALsbRsRVxkg98wQo3m3GSXelDwIAAAAAAAAAAADoLlESwHYGGSFVMdKJGQLwgscMk24i4sGAAAAAAAAAAAAAgC4RJQFspgqRxhFxbm4AbGCecVIVKS0MDgAAAAAAAAAAAGg7URLA+wa5EamKkXrmBcAOlmvbk2YGCQAAAAAAAAAAALSVKAngdeP8OjMjAPbgMeOkie1JAAAAAAAAAAAAQNuIkgD+W7UV6ToiLmxFAuCAbjNOmho6AAAAAAAAAAAA0AaiJIB/sxUJgCawPQkAAAAAAAAAAABoBVESULJqK9JVxki2IgHQJMuIuMtAaeZkAAAAAAAAAAAAgKYRJQElusgQ6dzpA9AC87XtSQAAAAAAAAAAAACNIEoCStHPEKnajHTi1AFooeVanPTgAAEAAAAAAAAAAIBjEiUBXTeIiOvcjtRz2gB0xG3GSVMHCgAAAAAAAAAAAByDKAnoqovcinTmhAHosPna9iQAAAAAAAAAAACAgxElAV3Sj4hxxkgnThaAgiwzTqq+Fg4eAAAAAAAAAAAA2DdREtAFgwyRqiCp50QBKNxtRFxHxEPpgwAAAAAAAAAAAAD2R5QEtNkwY6RLpwgAf3OfcdLUaAAAAAAAAAAAAIC6iZKANhrlQ9ZnTg8A3vWY3zcnRgUAAAAAAAAAAADURZQEtMk4H6o+cWoAsLEqTrrJOGlhfAAAAAAAAAAAAMAuRElA0/UzRroSIwFALZYZJ92IkwAAAAAAAAAAAIBtiZKApupniFR99ZwSANSuipPucgvhg/ECAAAAAAAAAAAAmxAlAU0zWNuMJEYCgMO4FScBAAAAAAAAAAAAmxAlAU0xyIehL50IABxNFSfdRMTMEQAAAAAAAAAAAABvESUBxyZGAoDmuc/vz1NnAwAAAAAAAAAAALzks6kAR1LFSJOI+L+CJABonLOI+GdGSSPHAwAAAAAAAAAAADwnSgIOTYwEAO0hTgIAAAAAAAAAAABe9Gm1WpkMcAhVjHQtRILGmUfE4o0P9ZBf+9CPiOEb/3+r//2pXzLQKPf5/XzqWAAAAAAAAAAAAKBsoiRg38RIsB+Pz2Kh54HA8/+5Co9mHTmLQX6te77BZfTs3z853MeDIoiTAAAAAAAAAAAAoHCiJGBfxEiwmeVaNLS+nWi2tslo9s5WI963vp3ptb+v/tozS/gQcRIAAAAAAAAAAAAUSpQE1E2MBH/3tNVofVvR0wP8QqPmeh4q9de2NFV/f1r6gGDNbX7/fzAUAAAAAAAAAAAAKIMoCahL9YD+VUR8NVEK9BQdzdbCo4XgqAj9tWDp+V9FS5RInAQAAAAAAAAAAACFECUBu3qKkaqvnmnSYfMMjKZrwdGDB+95x+DZ11OwdGZwdNxt3hsIMwEAAAAAAAAAAKCjREnALq5yG4IYia5YZmw0WwuQhEfsy1OwNHz21xMTpyOq31Nv8kucBAAAAAAAAAAAAB0jSgK2Mc4YyYPztNV6fPTwLESCJhitRUujDJcEoLTVU5x07QQBAAAAAAAAAACgO0RJwCZG+VDxqanRIvO1+GgqPqLF+hknDde2K505UFrkMcOkiUMDAAAAAAAAAACA9hMlAR8xzBjJw+803f3a1qOnL+i69UjJViXaoIpFrzIUBQAAAAAAAAAAAFpKlAS8ZZAbDS5NiQYSIMHrBmuxklCJprrPOMnv3wAAAAAAAAAAANBCoiTgJf18SPjKQ+w0xDwfWp8KkGBr65uUhrbf0SC3ec+xcCgAAAAAAAAAAADQHqIk4LlxRNyIkTii5Vp8NM0vYD9Gz7YpnZgzR7LM+48bcRIAAAAAAAAAAAC0gygJeDLKB4FPTYQDe1yLj2xBguMaPAuVfE/g0KrvCdcRMTF5AAAAAAAAAAAAaDZREjDIGOm8+ElwKPO1CGlqIwY0Wv9ZpHTmuDiQ+4yTbMsDAAAAAAAAAACAhhIlQbmqB82vIuKrXwPsmQgJumW09iVSYt9uM056MGkAAAAAAAAAAABoFlESlGmc25F6zp89eIyIOxESFONiLVI6dezswTLvW64NFwAAAAAAAAAAAJpDlARlGeUDvTZbUKflswjJNgsoVz+/1zyFSid+LVCjxwyrp4YKAAAAAAAAAAAAxydKgjL0c8PApfOmJvdrIdLMUIFXDJ5tUrKhjzrcZ5wkggUAAAAAAAAAAIAjEiVB913ldiQPgrOLx7UI6c4kgS2tb1E6NUR29C2j64VBAgAAAAAAAAAAwOGJkqC7Rvmgroe+2dbTNqQ72yiAPRg8i5TEs2zjMQNswSwAAAAAAAAAAAAcmCgJuqefMdKls2VDy7UIaWrzBHBgF2uR0onhs6EqpB2LaAEAAAAAAAAAAOBwREnQLeMMkmyb4KMeM0KaRMTM1ICGGGacdGHjHxtY5n3QtaEBAAAAAAAAAADA/omSoBuG+RDumfPkA+YZId3ZKAG0wGBti9K5A+MDHjPUnhoWAAAAAAAAAAAA7I8oCdqtHxFXEfHVOfIOIRLQBf21DUoCJd5zm/dJC5MCAAAAAAAAAACA+omSoL1GGZmcOENe8TMjpDsPZAMdJFDiI5YZJk1MCwAAAAAAAAAAAOolSoL26eeDtR7A5iVCJKBEAiXecx8RY9sCAQAAAAAAAAAAoD6iJGiX6mHam4joOTfWzDNUu/OwNYBAiTd9i4hrIwIAAAAAAAAAAIDdiZKgHQYZnZw5L5IQCeB9T4HSVUScmhdpnr8mpgYCAAAAAAAAAAAA2xMlQfNd54OztiPxmBFSFSPNip8GwGYGa4HSidkREd/zPmthGAAAAAAAAAAAALA5URI01zDjE5sdyrZcC5FsdACoR/U9dpxfot+yPeavA99jAQAAAAAAAAAAYEOiJGim6q39X51N0X6uxUgA7M9Ffl2acdFsTQIAAAAAAAAAAIANiZKgWWxHKlu1reEmY6SH0ocBcGD9jJOufB8ulq1JAAAAAAAAAAAAsAFREjSH7UhlWq5tRPIQNEAzDDNOqb56zqQ4tiYBAAAAAAAAAADAB4iS4PhsRyrTfG0rkoeeAZprnBuUzp1RUWxNAgAAAAAAAAAAgHeIkuC4bEcqy9NWpCpGmpU+DICWGaxtTzpxeMWwNQkAAAAAAAAAAABeIUqC47AdqSy2IgF0y0XGSbYnlcHWJAAAAAAAAAAAAHiBKAkO7yoi/jT3zrMVCaD7Bvl9vQpWes6782xNAgAAAAAAAAAAgDWiJDicQW5HOjPzTnvMEGnioWWAoozzy/f5bpvnOQuOAQAAAAAAAAAAKJ4oCQ5jnKGKLQrd9TPPeFr6IAAKN8ztSZelD6LjvuXWJAAAAAAAAAAAACiWKAn2q58bc87NuZOWeb5VjPRQ+jAA+C/9jJOqMPnEaDqp2pp04R4AAAAAAAAAAACAUomSYH9GEXFnO1InPeZ2hOp8F6UPA4B3jfPrzKg6Z5n3BDelDwIAAAAAAAAAAIDyiJKgfv18OPV3s+2c+zzbaemDAGArw9yedGl8nfMzwzOxMgAAAAAAAAAAAMUQJUG9qoeNJxFxaq6dcpsx0kPpgwCgFoMMWK5sVOyUamvShXgZAAAAAAAAAACAUoiSoD7Vg8V/mmdnVA8W3+SXrQcA7EN/LU46MeHO+J5nCgAAAAAAAAAAAJ0mSoLd9XM70rlZdsJjbkW6EyMBcEBPcZJti90wz61JtiwCAAAAAAAAAADQWaIk2M0o45WeObbePLciTUofBABHNco49swxtN4yQzP3FgAAAAAAAAAAAHSSKAm2Vz0w/NX8Wu8+z3Ja+iAAaJRRbk+6dCytd5txkg2MAAAAAAAAAAAAdIooCTY3yDfe22DQbmIkANpgkN+vxEntNs/IbFb6IAAAAAAAAAAAAOiOz84SNnKRD5MKktqr2lbwv7mBQpAEQNM9ZMzyS34Po51OI+Kv3JgEAAAAAAAAAAAAnWBTEnzcTUT8bl6tdZubJh5KHwQArTbIsKUKlXqOspV+5vktSh8EAAAAAAAAAAAA7SZKgvdVD//e5RvuaR8xEgBd1M846Uqc1EqPaxs4AQAAAAAAAAAAoJVESfC26mHRiYd9W0mMBEAJxEnt9iXvNQEAAAAAAAAAAKB1REnwuipo+Wo+rSNGAqBE4qT2us1zW5Q+CAAAAAAAAAAAANpFlAR/Vz3UexcRZ2bTKmIkAPj3fcxNRFyaRavMI2IcEbPSBwEAAAAAAAAAAEB7fHZW8F+GGbUIktrjZ0T8kg/yCpIAKN0ivyf+ksEu7XAaEdM8OwAAAAAAAAAAAGgFURL8x1VE/BURPTNphfuI+DUiLsRIAPA3D+Kk1qnuQX/kpisAAAAAAAAAAABovE+r1copUbp+Pvx5WfogWqKKka5zmwAA8DGDiJjYBtka84gY5eYrAAAAAAAAAAAAaCSbkijdMOMWQVLzPUbEb/mAriAJADbzkN9Df83Al2Y7zTMbOicAAAAAAAAAAACaSpREyS4ybjn1q6DRqhjpS254uCt9GACwo+lanPRomI3Wi4i/ImJc+iAAAAAAAAAAAABoJlESpbqOiH/kw5400zIivuWGgIkzAoBaTTP4/SJOarwf7oUAAAAAAAAAAABook+r1crBUJJ+PtR57tQb7XuGY4vSBwEAB1DdH13ll2C7uea55cr9EQAAAAAAAAAAAI0gSqIkTxt3Tp16Y/3MB6IfSh8EABxBFSfdRMSl4TfWMsOkWemDAAAAAAAAAAAA4Pg+OwMKUT28ORUkNdZ9RPwaEReCJAA4mmoDzzgifsnvzTRPtcnqrzwnAAAAAAAAAAAAOCpREiWoNu/8Mx/ipFkeI+LLWjQGABzfQ35v/jW/V9M8P3IDKAAAAAAAAAAAABzNp9VqZfp0WfWw5qUTbpxlRNzk16L0YQBAw1WB97XAu5Huc9Ok+ykAAAAAAAAAAAAOTpREV/Vz886pE26cn/lw80PpgwCAFulnmPS7Q2ucxwyTZqUPAgAAAAAAAAAAgMP6bN500DAfyhQkNcs8In7Nh2YFSQDQLouMin/J7Tw0x0nG+BfOBAAAAAAAAAAAgEMSJdE1F/lQ5omTbYxlRPyRsdi09GEAQMtVYfEoIn7LDT00Qy8i/pHhGAAAAAAAAAAAABzEp9VqZdJ0RfUQ5p9Os1Fu81wWpQ8CADqon9/nvzrcRqnuv8alDwEAAAAAAAAAAID9EyXRFZOIuHSajTHPh5RtRgKA7hvkvdiZs26M+9wgKgwHAAAAAAAAAABgbz4bLS1XvaF/JkhqjGVE/BERQ0ESABTjISJGEfFbRDw69kY4y3uxYemDAAAAAAAAAAAAYH9sSqLNhvlW/lOn2Ai3uR3JG/kBoFz9vB/46tdAIywzGJuVPggAAAAAAAAAAADqJ0qirZ428fSc4NFVGxHGNiMBAGsGGY+fGcrRLTMUmxQ+BwAAAAAAAAAAAGr22UBpobEgqRGqB1y/5UPHgiQAYN1Dbuj5kvcMHE91z/wjwyQAAAAAAAAAAACojU1JtE31MOWfTu3o7jMOeyh8DgDA+/oRcRMRl2Z1dLd5DwcAAAAAAAAAAAA7EyXRJhMPsx7dMsOwSeFzAAA2N8p7iBOzO6qfGSYtCp4BAAAAAAAAAAAANRAl0Qbert8MHmAFAHbVz8D5q0ke1TwjMfd1AAAAAAAAAAAAbE2URNNVD65OI+LUSR3NY8ZI00KvHwCo3zC3JrnHO5553uPNSh0AAAAAAAAAAAAAu/lsfjTYQJB0dN/zoWFBEgBQp1neY3wz1aM5zXu8YaHXDwAAAAAAAAAAwI5sSqKpnkKYnhM6CtuRAIBDGeTWpDMTP4pl3vfdFXjtAAAAAAAAAAAA7MCmJJpIkHRctiMBAIf0EBGjiPgjAxkOq7rn/keGSQAAAAAAAAAAAPBhNiXRNNXDkD+cylHYjgQAHJutScdVhWE3JQ8AAAAAAAAAAACAj7MpiSYRJB2P7UgAQBPYmnRcf2YUBgAAAAAAAAAAAO+yKYmmuMqHIDks25EAgKaqtibdRcSpEzq427xHBAAAAAAAAAAAgFfZlEQTTARJR2E7EgDQZA95r/LNKR3cZd6j9wu7bgAAAAAAAAAAADZgUxLHNsmHHjkc25EAgLYZ5n2jrUmHNY+IUUQsSrpoAAAAAAAAAAAAPsamJI5JkHR4P21HAgBaaJb3MN8d3kGd5n2jjUkAAAAAAAAAAAD8jU1JHEM/H270pvvDWeZ2pLtSLhgA6KxRxu0njvhgbEwCAAAAAAAAAADgb2xK4tAESYd3n5sFBEkAQBdM897mp9M8mNO1bVUAAAAAAAAAAADwL6IkDkmQdHjf8q32D6VdOADQadXGnouI+C03QrJ/J2tBGAAAAAAAAAAAAMSn1WplChyCIOmw5hExzjfaAwB02SAiJhFx5pQPYpnRu/tMAAAAAAAAAACAwtmUxCEMBEkHdetBUQCgIA957/PNoR9Ez8YkAAAAAAAAAAAAwqYkDmCYDy32DHvvlrkd6a7j1wkA8JpRbk06MaG9szEJAAAAAAAAAACgcKIk9kmQdDjziLjITQEAACXrZ5h07lfB3gmTAAAAAAAAAAAACvbZ4bMngqTD+Z7zFiQBAEQsMtb+wyz2rpf3/Bcdv04AAAAAAAAAAABeYFMS+yBIOoxlPgA6LeFiAQC2MMytSaeGt3dfctYAAAAAAAAAAAAUwqYk6iZIOoz7iBgIkgAA3jSLiFFE3BrT3v2IiHHHrxEAAAAAAAAAAIA1oiTqJEg6jG/5cO2ihIsFANjRImOZL7lpkv0RJgEAAAAAAAAAABTk02q1ct7UQZC0f9VDtBe2IwEAbK26Z72LiBMj3KsqAJt0+PoAAAAAAAAAAACKFzYlURNB0v7N1+YMAMB2ZnlP9dP89srGJAAAAAAAAAAAgAKIktiVIGn/vuecH7p+oQAAB7DI7ZN/GPZeCZMAAAAAAAAAAAA67tNqtXLGbEuQtF/LiLiKiEmXLxIA4Ijcz+7fF/ezAAAAAAAAAAAA3WRTEtvyAOd+zSNi5AFOAIC9mkXEICLujXlvbEwCAAAAAAAAAADoKFES2xAk7dfPDJJmXb5IAICGWOS913cHsjc3+TMEAAAAAAAAAAAAHSJKYlOCpP36FhEX+XAsAACHcxURXyJiaea16+XPEMIkAAAAAAAAAACADvm0Wq2cJx8lSNqf6uHXcUTcdfUCAQBaYpj3ZCcOrHZLG0EBAAAAAAAAAAC6w6YkPqofERNB0l7M8+FMQRIAwPHNMky6dxa1szEJAAAAAAAAAACgQ0RJfEQ/Hx48Na3a/fS2eACAxlnkPdp3R1M7YRIAAAAAAAAAAEBHiJJ4jyBpf75FxEU+9AoAQPNcRcQX51I7YRIAAAAAAAAAAEAHfFqtVs6R1wiS9mOZD7hOunhxAAAdNMz74p7DrdVjzlakDwAAAAAAAAAA0EKiJN4yEyTV7jG3I806dl0AAF0n2N+PeUSMhEkAAAAAAAAAAADt89mZ8YqJBy5rN883wQuSAADaZ5HxzK2zq9Vpxl79Dl0TAAAAAAAAAABAEURJvKQKki5Npla3GSR5AzwAQHtV93LjiPjmDGslTAIAAAAAAAAAAGghURLPCZLq90c+vAoAQDdcR8SXiFg6z9qc5s8iAAAAAAAAAAAAtMSn1WrlrHhyFRF/mkZtljlTD1cCAHTTMDf89JxvbW4F/QAAAAAAAAAAAO0gSuJJ9eDfD9OoTRUkjSJi1pHrAQDgZYOIuMtNP9RDmAQAAAAAAAAAANACnx0SgqTazfOt+YIkAIDue8gY/d5Z1+YyN44CAAAAAAAAAADQYDYlUcUzfxU/hfpUD6NeRMSiKxcEAMCHTTKooR5fcqYAAAAAAAAAAAA0kE1JZauCpGnpQ6jRbb4lX5AEAFCmagPpH86+Nj8y+AcAAAAAAAAAAKCBbEoq1yAiZhHRK30QNfkWEdeduBIAAHY1zqCG3S0z/J+ZJQAAAAAAAAAAQLOIksrUzw1Jp6UPoiZfImLSiSsBAKAuVUhz5yUAtRAmAQAAAAAAAAAANJAoqTyCpPos8y34d125IAAAajXMe29h0u4ec56Ltl8IAAAAAAAAAABAV3x2ksW5ESTVYrn29nsAAHhJtdlnEBFz09nZSQZe/ZZfBwAAAAAAAAAAQGeIksoyiYjL0odQg3kGSbPWXwkAAPu2yHtHYdLuTvNnGgAAAAAAAAAAABpAlFSOsSCpFoIkAAA29RQm3Zrczs6FSQAAAAAAAAAAAM0gSipDFST9KH0INXgKkhatvxIAAA5tkfflwqTdVS9buGr7RUBhhvnzNAAAAAAAAAAAHfJptVo5z26rHvyZRkSv9EHs6DYfIgUAgF1NbDGtxRdbk6AxRvk1WPs6eefDLXML8SL/Oss/v/AiEAAAAAAAAACAlhAlddsgH+oRJO1GkAQAQN1sM93dMiOIWdsvBFqoegHKRX6d1vzxHyPiLgOlO784AAAAAAAAAACaS5TUXf18gKfuh4NKI0gCAGBfhEm7W2Yc8dD2C4EWGOTvW+MPbEGqyzLDpBsBIgAAAAAAAABA84iSuqsKks5KH8KOvkTEpNVXAABA0wmTdjfPjUmLtl8INFT139dVRJwf+ePNM07yczoAAAAAAAAAQEOIkrqpekDnsvQh7EiQBADAoYxyE0jPxLd2n3ME6lP9N3XdwBeePObn8jM7AAAAAAAAAMCRiZK6x5vWdydIAgDg0Ia57VSYtL3b/HkI2M0gNxIdezPSe+a5wWna7I8JAAAAAAAAANBdn51tp4wESTsTJAEAcAyzvJ9fmv7WLkVJsLOr/P2o6UFS5TQi/pkBVb8BnwcAAAAAAAAAoDg2JXWHN6vvpnr488IblgEAODL39bv71X09bGyQL+g4a+noHjNK9N8+AAAAAAAAAMAB2ZTUDf18eMiDi9tZ5lvpPbwEAMCx2Zi0u7uMu4CPucjfe9oaJFVOcmvSdQM+CwAAAAAAAABAMURJ3VA9dHda+hC29BQkzVr56QEA6CJh0m56+dKGfpsvAg7kKiL+0aGXnHz13z8AAAAAAAAAwOF8Wq1Wxt1u1cM2l6UPYUuCJAAAmqyf2zy9gGA793m/D7ysy3+eMM///hcN+CwAAAAAAAAAAJ1lU1K7jQVJWxMkAQDQdIu8Z507qa2cRcRNCz83HELXX3BymlGnjUkAAAAAAAAAAHtkU1J7DSPir9KHsCVBEgAAbWJj0m6+ZIAB/FtJG5dtTAIAAAAAAAAA2CNRUjtVDyU+RESv9EFsQZAEAEAbCZN2879+BoB/KSlIeiJMAgAAAAAAAADYk88G20pTQdJWBEkAALTVIu9l505wK9MMu6BkVwUGSZExp21pAAAAAAAAAAB7IEpqn4m3o29FkIaIMZoAACAASURBVAQAQNsJk7bXyzAJSnUREX8WfP3nEXHTgM8BAAAAAAAAANApn1arlRNtj3FE/Ch9CFsQJAEA0CX9DGy8rGBzt/lzFZRkkD8P27gc8VtE3DXgcwAAAAAAAAAAdIIoqT2GEfFX6UPYgiAJAIAuEiZt70tuoIVSVL9XnDntf1lmpLVowGcBAAAAAAAAAGi9z46wFZ4eOGQzgiQAALqqeqD+Iu952cxNvvQBSnAlSPovPZuSAAAAAAAAAADqY1NSO8y8AX1jgiQAAEowzBcY9Jz2Rh5zdral0GWD/JnY7w9/95s4CQAAAAAAAABgdzYlNd+NIGljgiQAAEoxy3tfG5M2cyJIoAA3gqRX3eRWagAAAAAAAAAAdiBKarZxRPxe+hC2cCVIAgCgIMKk7ZxFxHUbPzh8QPV7wrlBveok/+wAAAAAAAAAAIAdfFqtVubXTMOImHqr8ca+RMSkZZ8ZAADq4GeI7fyac4MumWZ4x+uqkHMQEQszAgAAAAAAAADYjk1JzdTPsMbDhJsRJAEAUDIbk7Zzl2ECdMVIkPQhPduSAAAAAAAAAAB2I0pqppuIOC19CBsSJAEAwL/DpLE5bKSXYRJ0hdDm467yxTAAAAAAAAAAAGxBlNQ81QOEl6UPYUN/CJIAAOD/u8ton487zZdDQNtVW7/OneKHVVHiRUs+KwAAAAAAAABA44iSmmUYET9KH8KGbj08CAAAfzMRJm3sd3ECHWBL0ubMDAAAAAAAAABgS59Wq5XZNUM/ImYRcVL6IDZwm5ulAACAl429+GAjy3xZxEOLPjOse/DnClv5xX/3AAAAAAAAAACbsympOSYeHNqIIAkAAN43yXtnPqYXEXdmRUsN/bnC1mxJAwAAAAAAAADYgiipGa4i4rz0IWxgnjMDAADeNxYmbeQ0Im5a9HnhiRd3bM/sAAAAAAAAAAC28Gm1WpnbcVVvMp7mG7l5XxUkjSJiYVYAALCROy9D2MhvtibRMrOM6tjO//FnDQAAAAAAAAAAm7Ep6bj6ETERJH3YoyAJAAC2Ns7In4+pflYbmBUt0Rck7WzU8s8PAAAAAAAAAHBwoqTjuvHQ0IctI+JCkAQAAFtb5EP3wqSP6dmURIsMHdbOzBAAAAAAAAAAYEOipOOpApvLUi9+Q8t8eHLWqk8NAADNs8ifRZbO5kOql0hct+Bzgi0/uzNDAAAAAAAAAIANiZKOYxARkxIvfEtXgiQAAKjNQz58L0z6mK9iBVrAlp/dmSEAAAAAAAAAwIZEScdxFxG9Ei98C18EXAAAULtZbkziY6qfSfpmRYP59bk7f04DAAAAAAAAALAhUdLhXUfEaWkXvaXvgiQAANibab4EgPed+NmEhjtzQLWwFQ0AAAAAAAAAYAOipMOqHm75WtIF7+A2Iq5a++kBAKAdqtDmm7P6kHM/owAAAAAAAAAAAPzHp9VqZRyH0Y+IWb5hm7fNM+BamBMAABxEFSddGvW7lhExjIiHhn9OyuMPd+rxa26RAwAAAAAAAADgA2xKOpyJIOlDBEkAAHB447wX5229iLgzIxpm6EBqM+rIdQAAAAAAAAAAHIQo6TAuIuK8hAvd0TIfhhQkAQDA4Y2ESR9yGhHXLficlKPvrAEAAAAAAAAAOAZR0v4NcksS76segpyZEwAAHMUiXxKwNP53fbVRBQAAAAAAAAAAKJ0oaf+qIKnX9YuswRdBEgAAHN1MbPNhExtqAAAAAAAAAACAkomS9usqIs66fIE1+W6bFAAANMYsXxrA204i4tqMAAAAAAAAAACAUomS9mcYEX929eJq9DPjLQAAoDkm+fIA3vZ7RFyYEQAAAAAAAAAAUCJR0v7Y/PO+eUSMm/4hAQCgUFf5EgHeVv3s1zcjAAAAAAAAAACgNKKk/biOiNMuXliNlvlG8UVnrggAALpnnC8T4HU9L6UAAAAAAAAAAABKJEqq3zAivnbtovZgFBEPnbsqAADolkW+TGDpXN90nnMCAAAAAAAAAAAohiipft6Q/b4vETFr+ocEAAD+5UFw8yHVz4L9FnxOAAAAAAAAAACAWoiS6nUdEadduqA9uBVuAQBA60zz5QK8rudnHQAAAAAAAAAAoCSipPoMI+JrVy5mT+4jYtzJKwMAgO6b5EsGeN25rVIAAAAAAAAAAEApREn18Ubstz16OA8AAFqvesnA3DG+qfrZsN/gzwcAAAAAAAAAAFALUVI9riPitAsXsifLDJIWnbw6AAAoyyjv8XlZz0srAAAAAAAAAACAEoiSdjeMiK9tv4g9u4qIWaevEAAAyrHIMInXndsUCwAAAAAAAAAAdJ0oaXfegP22WzMCAIDOqV468MWxvqn6Oajf4M8HAAAAAAAAAACwE1HSbq4j4rTNF7Bn84gYd/oKAQCgXJN8CQEv63lBAwAAAAAAAAAA0GWipO0NI+JrWz/8ASwjYtT5qwQAgLJd5csIeNl5RFyYDQAAAAAAAAAA0EWipO3dtPWDH0j14N2iiCsFAIByLfLef+nXwKuqnx37Df1sAAAAAAAAAAAAWxMlbad6G/hZGz/4gfwREdMirhQAAHiIiHHxU3jdSURcN/XDAQAAAAAAAAAAbEuUtLmBB8re9NMWKQAAKM5dRHx37K/6PSJGDf1sAAAAAAAAAAAAWxElbW4SEb22fegDefSGdAAAKFa1Ufbe8b9q0tDPBQAAAAAAAAAAsBVR0mYuIuKsTR/4wKr5LIq6YgAAYF31M8HSRF50YusuAAAAAAAAAADQJaKkj+t7s/Wb/oiIWYM/HwAAsH+LDJN42deIGJgNAAAAAAAAAADQBaKkj6veaN1ry4c9sJ8RcVPUFQMAAK+ZRsQ303mVl10AAAAAAAAAAACdIEr6mFFE/N6GD3oEjxExLu6qAQCAt1Qvdbg3oRed+RkKAAAAgP/H3t1ftZFkfQC+O2f+l94IYCKAjQBtBLARwERgJgLjCKyJwDiCwREYIhiIYCCClSKY97RdGgsMmI9udXXf5zmHw36872ypSkjV3fdXFwAAAADGQCjpaXQBethBRCxqHRwAANCb5lphafrv1VxjTiscFwAAAAAAAAAAwJMJJf3YcUTs1D7InvwWEZcpXzkAAPAjixJM4nsTh18AAAAAAAAAAABDJ5T0uO2IOKl5gD36pIgOAAD4gfOI+N0k3eswImYVjgsAAAAAAAAAAOBJhJIeNy8nWHPbMiKOzAkAAPAETffZKxN1Lwc9AAAAAAAAAAAAgyWU9LDmxOr9WgfXs4OIWKSeAQAA4DkOyuEG3LZTQlsAAAAAAAAAAACDI5T0sNNaB9azdxFxnnoGAACA57oWvnnQSURMKx0bAAAAAAAAAADAg4SS7tcUhW3VOLCeXZW5AQAAeK7m4IdPZu07k4iYVzYmAAAAAAAAAACAHxJK+t62E7zvtYyIgwrHBQAADMdRRNxYr+8cRsSssjEBAAAAAAAAAAA8Sijpe/NyUjW3NR2Srs0JAADwCosSTOJ7uiUBAAAAAAAAAACDIpR0W3My9X5NA6rEJwVyAABAS84j4p3J/M6Orr0AAAAAAAAAAMCQCCXdJnjzvaWTzAEAgJY1nVivTOp3mnmZVjYmAAAAAAAAAACAewklfXNcTqbmtiaQtDAnAABAy47KIQh8MynBJAAAAAAAAAAAgOoJJX01Vfh1r98j4qzCcQEAAMN36TrsXm8iYrfCcQEAAAAAAAAAANwilPTVSTmRmm9uFAgCAAAdm0fEhUn+zryy8QAAAAAAAAAAAHxHKCliu5xEzW1HEbEwJwAAQMeaa4+lSb5lLyIOKhoPAAAAAAAAAADAd4SSIk4rGENtfo+I8+yTAAAAbMS1Lq330i0JAAAAAAAAAACoWvZQ0qycQM03VxFxbD4AAIANagI4n0z4LVvCWgAAAAAAAAAAQM2yh5J0SfreUW0DAgAAUmiuRZaW+pbmwIhpReMBAAAAAAAAAAD4R+ZQ0nE5eZpv3kXEpfkAAAB6sHBIwncmuiUBAAAAAAAAAAC1yhpKmirs+s6VOQEAAHp2FhGfLMItbyJiu6LxAAAAAAAAAAAAfJE1lHRcTpzmGyeSAwAANWiuTZZW4pbTisYCAAAAAAAAAADwRcZQUnPC9NsKxlGT3yPiMvskAAAAVVjo4vqdvYiYVTYmAAAAAAAAAAAguYyhJMVtt92YEwAAoDLziLiwKLe4bgMAAAAAAAAAAKqSLZS0GxGHFYyjJkflJHIAAIDarlWWFYyjFntlTgAAAAAAAAAAAKqQLZQ0r2AMNfk9Is6zTwIAAFCla92BvmM+AAAAAAAAAACAamQKJc3KydJ8tVTQBgAAVK45WOLKIv1jKyKOKxkLAAAAAAAAAACQXKZQki5Jtx1FxKKmAQEAANzjyKTc0hwuMa1oPAAAAAAAAAAAQFJZQklNEdtOBeOoxaeIOMs+CQAAwCBcRsQ7S/WPiW5JAAAAAAAAAABADbKEkk4qGEMtlgrYAACAgWk6395YtH8c65YEAAAAAAAAAAD0LUMoqemStFXBOGrRBLSus08CAAAwKItybcdXE4dvAAAAAAAAAAAAfRt7KGmqUOuWq3LCOAAAwNCcR8Qnq/aPNxGxXclYAAAAAAAAAACAhMYeSjrWJekWJ4sDAABD1lzTLK3gPxzCAQAAAAAAAAAA9GbMoaRpCSXx1e8RcWkuAACAAVsI4txyqFsSAAAAAAAAAADQlzGHkppA0qSCcdRgqXAPAAAYiXlEXFjMf7jWAwAAAAAAAAAAejHWUJIuSbcdlRPFAQAAxsD13je6JQEAAAAAAAAAAL0YayhJl6RvmhPEz2oZDAAAQAsuI+J3E/kP3ZIAAAAAAAAAAICNG2MoSZek245qGgwAAEBLmiDO0mR+0XRLmlUwDgAAAAAAAAAAIJExhpJ0SfrmXURc1zIYAACAFi0cSHGLbkkAAAAAAAAAAMBGjS2UpEvSN82J4fNaBgMAANCB04i4MLFf7OmWBAAAAAAAAAAAbNLYQkm6JH1zXE4OBwAAGDMdgr4xFwAAAAAAAAAAwMaMKZSkS9I3F+XEcAAAgLE7j4iPVvkL3ZIAAAAAAAAAAICNGVMoSZekb4SzAACATJproKUV/0K3JAAAAAAAAAAAYCPGEkrSJemb5oTwy1oGAwAAsAGLiJib6C+abkm7FYwDAAAAAAAAAAAYubGEknRJ+mopnAUAACTVdAi6sfhfuC4EAAAAAAAAAAA6N4ZQki5J38zLCeEAAAAZuTb86jAitmsYCAAAAAAAAAAAMF5jCCXpkvTVTTkZHAAAIKuziLiw+l+4PgQAAAAAAAAAADo19FCSLknfmAcAAADXRiu6JQEAAAAAAAAAAJ0aeijpSJekLy7KieAAAADZXUbEx+yTUOiWBAAAAAAAAAAAdGbooSQnYH+l0AwAAOCb5lpxaT50SwIAAAAAAAAAALoz5FBS0yVpq4Jx9K05Afw89xQAAADcsoiIuSn5wmEeAAAAAAAAAABAJ4YcStId6CvzAAAA8L0mlHRjXr4c6DGtYBwAAAAAAAAAAMDIDDWUpEvSV+8i4rqGgQAAAFRm4RCHLya6JQEAAAAAAAAAAF0Ycigpu2U5+RsAAID7neqW9MWxbkkAAAAAAAAAAEDbhhhKmkXEXgXj6Nu8nPwNAADAwxxq8bVb0kEF4wAAAAAAAAAAAEZkiKGkkwrG0LcbXZIAAACe5DwiLkyVa2kAAAAAAAAAAKBdQwslbeuS9MWJLkkAAABPJpATsaVrFAAAAAAAAAAA0KahhZIUkn3tknRawTgAAACGQrekr4SSAAAAAAAAAACA1gwplNR0STqsYBx9E8wCAAB4PoGcr52HZxWMAwAAAAAAAAAAGIEhhZIUkEVc6ZIEAADwItcR8dHUxXEFYwAAAAAAAAAAAEbg54G8hKnCqS/MAQAAwMud6MAb+6UT8XUFYwHGY7fcv2vbtc8rAAAAAAAAAKjXUEJJBxExqWAcfbqIiPO8Lx8AAODVVt2SsgeTTnQjBl7hoISQZuX3Ju7ZXZXP8PPyc2kBAQAAAAAAAKB///r777+HsAxN0cFWBePo03+EkgAAAF6t6RL0V/JpXJZ5WFQwFl6vCYZ8No+teFdCe9w2LUGkg9JtrQbN59jZ2g8AAAAAAAAA0IOfBjDpM4EkXZIAAABasuqWlNlEpyTgCZrw4mn53PxQUSApyudY0/XujzK+kxKeAgAAAAAAAAA2aAidkpowzl4F4+iTLkkAAADt0S0p4qbMA8OnU1J7dEr6arvMw2ENg3mGpnvSvPzoBAf0Zbb2vzu7M4a7/z46fPbRfCZe3vnPFnf+s7v/3jMIAAAAAAAAnq32UJJCsa9dku57WAkAAMDLnQ6w4L5t/42Is3G9pJSEktqTPZQ0La//TQVjeY2mEP+4fM4DtGW3fE6ufm+vBbzHdqjaeqDpsoSXru/8AAAAAAAAwBe1h5IUiemSBAAA0AWHYDgEYyyEktqTOZQ0K/fhtioYS1uaz7ijUDwPPN1sLWy0HkKamMPv3NwJKV2u/QYAAAAAACCRnyt+qc0Dv4MKxtGnC4EkAACATjRFkx+TH4SxV4puFexDbvMRdEe6z14pjj/SFQ5Yswoa7a6FjwSPnm+r/NzXJWoVWDpfCy15zgEAAAAAADBSNYeSjjwITHs6LwAAwCac6M77ZQ6OKhgHsHnTEta5r6B8LJp7i38k74IFma2HjlY/Y+oIV6uHAktXa92UzsvvRfbJAgAAAAAAGLp//f3337W+hOvkDwibLkmzCsYBAAAwZqfJg0nLUrCrIHS4mnsHn7NPQksyBVempSB8p4KxbMpHIUwYtVUHpNna7+yHng3BzZ2Qko5KAAAAAAAAA1Nrp6SZEwud3goAALAB2bslTUqR/ryCsQCbkTGQFGuf9YJJMA7b5TnCKoSU7TNtLFZdlfbXXs/FWkDpXHgeAAAAAACgbrWGko4rGEOfLpwICAAAsBHXpXtG5mDSsVASpJE1kLQimATDtR5CcqjZuO2VnzflVV6tBZSElAAAAAAAACrzr7///ru2MTUPF/+qYBx9+o9QEgAAwMa4DnUdOmRNYfbn7JPQkncj71ydPZC07qNgElRvuhZAOhBCYs0qpHRm/woAAAAAANC/nypcg+wFAbokAQAAbNaqW1Jm2TsWQwanAkn/OHQPEqq0W/Ykzf3x/0XEH6VbjkAS63bK++Jz6Zp0Vj7Tt80SAAAAAADA5tXYKek6+UPGX0uRCAAAAJujW1LEL+WanGHRKak9Y+6U1BT5v69gHLX5d0RcZp8E6NmBbki0aNVF6dTnOwAAAAAAwGbU1inpKPmDxxuBJAAAgF40YZxPyade1xAYp12BpAe5Dwf9OCh/fwvdkGjZqovSn2V/Py+hNwAAAAAAADpSYygps7GexgsAADAE8+SrlP2aHMYq+2fbY3bcj4ONuRtEOoyIiemnQ1sloPS5vO9OBZQAAAAAAADaV1MoaTsi9ioYR190SQIAAOjXeURcJF6DrVIwDIzHUfL7bU/xttyXBNoniEQtJuX993mtg9Ku1QEAAAAAAHi9mkJJxxWMoU8CSQAAAP3L3jFDtyQYj6kuSU+W/bMf2rRbPnsEkajVqoPSnyWgdCycCgAAAAAA8HI1hZIyFz4tFYkAAABU4bx0ss1qX1EmjMaxIMCTHeqYAa8yLZ85lyXo8cbnDwPRBJTeR8Rf5TpAQB8AAAAAAOCZagklHSR/SLk6ORIAAID+Ze+YoRgTxiF7V/LnMl/wfLOIOI2I/5Vgx445ZMD2IuJDeVYzF1YFAAAAAAB4mlpCSdkLnk4rGAMAAABfnSbvlpT9Gh3G4EiXkmc71CkOnmTVFek6Ij6Xvx0Yk0np9vWn7kkAAAAAAAA/VkMoqXnYv1/BOPrysTzABQAAoB6ZD4/YKp0PgOHS9edlFJ7Dw3bvdEXaMlcksN496UR4FQAAAAAA4Hs1hJKyP+w/qWAMAAAA3DaPiGXiOcl+rQ5D1hRM71jBF/HZB987Kt1i/tQVicSa7klvI+KvEs4T4AcAAAAAACiEkvp1oUsSAABAlZrT0M8SL01TdDytYBzA8x2YsxfbKt1gILtp6bh2XbrE7GWfEFjT7JM/R8SlMCsAAAAAAED/oaRZediflS5JAAAA9cp+zSbYAMPkb/d1dL8gs2nZ/zRhpPfJ793Dj+yU0N51CScJ9AMAAAAAACn1HUrKfIrcTUScVzAOAAAA7tcUGH5KPDfHFYwBeD4dTV5HqIuMtiPiNCL+FxFvI2LiXQBPtrUWTjoRTgIAAAAAALLpM5Q0Tf6QP/uJ2wAAAEMwT7xKO6VIGRgOXX5eb3foLwCeYRVG+isiDk0cvMqkhPqEkwAAAAAAgFT6DCUdJD5xcRkRZxWMAwAAgMc1HW6vEs+RbkkwLAI1rzcRyCQBYSTojnASAAAAAACQSp+hpKPEb7Xmge+ignEAAADwY5m7JWXucAxDJEzTDvPIWAkjweYIJwEAAAAAACn0FUpqHn7uJX6LZS5oAwAAGJrT0vE2oy3BJBgUnZLaMRvDi4A1wkjQH+EkAAAAAABg1PoKJWUuaPpUHj4BAAAwHKeJ10ooCQCGaVpCEMJI0L/1cNKR9QAAAAAAAMair1DSceJ3kC5JAAAAw5P5Wu7Aie4wGDolASsnJfzw1oxAVZpw0gfhJAAAAAAAYCz6CCU1xRFbSd9BNxFxXsE4AAAAeJ7r0vk2o4luSTAYE0vVitkIXgN5Ha2FkXwmQL22Sjjp3PcOAAAAAAAwZH2EkjKf/KZLEgAAwHBl75YEANRrVsINHxIfCgZDtBcRnyPiNCK2rSAAAAAAADA0QkmbsywPlQAAABim89IBN6N9RZIAUKVpue/8uYQbgGE6jIjLiDgpf9cAAAAAAACDsOlQUnOy8iTpW+MsIhYVjAMAAICX0y0JAKjFcURclzADMHzN87O3JZxk7w0AAAAAAAxCH6GkrDIXrgEAAIxF5g64WTsfA0BtZiW08D7xIWAwZlsR8Ufp1KpbKQAAAAAAUDWhpM24Kg+JAQAAGLamA+7HpGu4oygSAHo1LQHpz+V7GRi3vfJs6cQ6AwAAAAAAtdpkKOkg8amNuiQBAACMR+ZuSZk7IANAn5qOhdcRcWgVIJXmudrb8vc/s/QAAAAAAEBtNh1KymgZEWfe+QAAAKNxHhE3SZfzqIIxAEAm22Xv8SHxoV9AxFbpkjYvXdMAAAAAAACqsKlQ0jRxKKkJJC0qGAcAAADtydoRd6cURwMA3TuOiMuI2DPXQPGmfC7oYAoAAAAAAFRhU6Gkg8SnOGYtVAMAABiz08Sre1zBGABgzFbdkd7rjgTco+ma9Ec5FE/XJAAAAAAAoFebDCVldFNOrAMAAGBcmo64H5OuqVPZAaA7uiMBT7UfEdf25wAAAAAAQJ82EUqalgcjGemSBAAAMF5nSde2OZl9t4JxAMCY6I4EvMSkdE2a65oEAAAAAAD0YROhpMwntJ1WMAYAAAC6cVY65GZ05D0FAK050B0JeKU35XNkZiIBAAAAAIBNEkrqzqeIWIz1xQEAAPBF1m5Jih0B4PWmZS/xh+5IQAuajqafI+LEZAIAAAAAAJuyiVDSftLV1CUJAABg/OZJ13gnIrYrGAcADNVu6WqS9f450J235fPFfh0AAAAAAOhc16GkrF2SlolPywYAAMjkOiKukq541mt+AHitpovJn6WrCUAXdkowyZ4dAAAAAADolFBSN3RJAgAAyCNrt6SjCsYAAEMyjYjz0sUEoGuTiPgj8fUKAAAAAACwAUJJ3RBKAgAAyCNrp9zm9PXtCsYBAEOwWzos7lktYMPelK5J9u4AAAAAAEDrugwlHZRT2LK5Kg93AAAAyGERER+TrnXWw0gA4DmOI+LPpPfLgTrslGdX9u8AAAAAAECrug4lZaRLEgAAQD5ZuyUpagSAh03L/eL35gioQBOM/CMiTiwGAAAAAADQli5DSbOkq5S1EA0AACCz5lpwmfD175WCawDgtt2IOI+IQ/MCVOZt+XyyjwcAAAAAAF6tq1BS88B1K+HyXETEdQXjAAAAYPOyds7VLQkAbpuVgv8d8wJUqjlc4LI8zwMAAAAAAHixrkJJR0mXJGsBGgAAAEJJAEDEcUR8joiJuQAqt1UClPbzAAAAAADAi3UVSpolXZKzCsYAAABAP5qTxm8Szv1+BWMAgBo0AeX3VgIYkCZA+UcJVAIAAAAAADxbF6Gk7YjYSbgUnyJiUcE4AAAA6E/Wwyqcrg5AZtMSTj70LgAG6n3izq8AAAAAAMArdBFKylqIpEsSAAAAWQv5hJIAyGo3Is6THtQFjMthCVhOrSsAAAAAAPBUXYSSZglnf+kEOQAAAEoR31XCich4LwAABJKAsdkpn2vbVhYAAAAAAHiKtkNJzelp+wlnXpckAAAAVjIeWrFVCrMBIIujUrg/seLAyOyUwxbs7wEAAAAAgB9qO5SU9WRkoSQAAABWsl4j6pYEQBZNIOmDQBIwYpMSvLTHBwAAAAAAHtV2KOkg4XQvhZIAAABYcx0RVwkn5KiCMQBA105KIAlg7Jpg0mf7fAAAAAAA4DE6Jb2eQBIAAAB3nSackZ2ImFYwDgDoSvP9/tbsAsl8EEwCAAAAAAAe0mYoaTcithLOtFASAAAAd2W9VszYQRmAHJpA0qG1BpL6UDrFAQAAAAAA3NJmKCljl6SlUBIAAAD3uI6Iq4QTk/HeAADjJ5AE8LVTXMaOsAAAAAAAwCPaDCVlPA1ZIAkAAICHZLxmFEoCYEymAkkAtxwKJgEAAAAAAOvaCiU1D2f3Es7seQVjAAAAoE4ZQ0lbEbFbwTgA4LWm5f6vQBLAbYJJAAAAAADAP9oKJWU9CVmnJAAAAB5yGRE3CWdHtyQAhm4VSNqxkgD3EkwCAAAAAAC+EEp6uU8RsRjq4AEAANiIjIdZHFQwBgB4KYEkgKcRTAIAAAAARGhKHAAAIABJREFUAFoLJWUsONIlCQAAgB/JWKS3V8EYAOAlBJIAnkcwCQAAAAAAkmsjlLQdEVsJp1EoCQAAgB+5jIhlwlnSLQmAIZoLJAE8m2ASAAAAAAAk1kYoaZZw+q4iYlHBOAAAAKhfxkMtMt4rAGDYTkthPQDPJ5gEAAAAAABJCSW9jAcrAAAAPJVQEgDUTSAJ4PUOS8c5AAAAAAAgkZ9beKkHCd8w5xWMAQAAgGHIGEraiYipLsMADIBAEjW6euI+ajsitqwgFXkTEZcO9wMAAAAAgDxeG0rajYhJsvfLTXmgAgAAAE/1KSL2k83WLGkgC4DhOBFIomMX5R9/XX6iPF9YBY4WHT1v2C0B8Si/d8u/3i4/0xIihy58KP9MwSQAAAAAAEjgtaGkWcI3iYIqAAAAnussYSjpwDU0ABU7ioi3FohXWpZQ0SpodF7+cec9T+zdoNNDe7LpWoBpdy20tLeBMTJugkkAAAAAAJCEUNLz9f0wEQAAgOHJeC2Z8Z4BAMNwtFYwD091tRZAurzT8Wio1oNUd4NLq4DSbC2wpLsSzzFf+1sBAAAAAABGSijpeZZOeQYAAOAFrksha6ZCzq1SvHpdwVgAYGW3FMrDY25KWGcVqMgYML8uP3df+2wtqNT8nvQ0Puo3Ke+fmWASAAAAAACM12tCSbsJHzbpkgQAAMBLnSc8Xb4pQDytYBwAEOWe9rkQBfe4KQeSrYJIQtUPO7/zrGR7Lag0K8F0WJmUv63dEXQWAwAAAAAA7vHTKyYlW5ek0CUJAACAV8h4TZnx3gEAdZqWoKxAEo1lRHyKiF8j4pcSrDku+zWBpOe5Ln9bR2Ue/x0Rv5X5hShBtfPyOQwAAAAAAIzMazolZSws0ikJAACAlzovBbCZiqGFkgCoRcaOhdy26oZ05l5/py7Lz7yEUJr94EH5EQrMa6e8J46yTwQAAAAAAIyNUNLTXTkhEQAAgFdqCmD3E03iVjkx3/U0AH06FUhKaxVEOi1BGTZrsRYEizsBpS1rkc5heU8cZ58IAAAAAAAYk59e+Fp2E55o5+REAAAAXuss4QzuVjAGAPI6LoXw5NEEkX6PiH+XcPSxQFI1zst6NOvy34j4WDqJkscb3ZIAAAAAAGBcXhpKytYlKYSSAAAAaEHGa8uM9xAAqEPzHfTeWqSwLAGX/wgiDcZZCadMI+LXiPiUfUISmTu4AAAAAAAAxkMo6ekynmYNAABAu67L6f2ZCCUB0Idd93RTuCqBlu0ScHG42DCdRsRBRPwSEe8S7pezmZS/1Wn2iQAAAAAAgDF4aSgp2wlmFxWMAQAAgHHIViC9o+AQgA2blpDDxMSP1qor0m5Z60X2CRmJJsB/UkJm//VsZtQmQoQAAAAAADAOLwklNQ+DtpKtvxM1AQAAaEvG4jvdkgDYpNMSimVclqWLzi+6IqVwVvaQv5QQGuOzUz6vAQAAAACAAXtJKCljIZGHmwAAALQl4zVmto7LAPTnOCL2zf+o3ETEr+XAtJPSTYc8rksI7f9KKG1p7UflsKwvAAAAAAAwUC8JJWUrJGoecF1WMA4AAADGYRERV8nWUqckADah+b55b6ZHYz2MdFr2UOS1KKG0beGk0Zk7xAAAAAAAAIZLp6Qf0yUJAACAtp0lm9G9CsYAwLhNE36/jtXdMBKsE04an0n5W59mnwgAAAAAABiil4SSdpKttFASAAAAbct4ren0cwC6dFYK2xkuYSSeQzhpXHb83QMAAAAAwDA9N5SUrUtSCCUBAADQgYzXmhnvKQCwGSe68g3aUhiJVxBOGo/9iDjOPgkAAAAAADA0QkmPax5eXdY8QAAAAAbrItnS6ZQEQBeae9ZvzewgLUuIRBiJNqzCSc2e86MZHawT1w0AAAAAADAszw0lZXsQoEsSAAAAXcl2zalTEgBtmwqzDNbH8rzhpIRJoC3XEXEUEf9OeAjAGEzK5/o0+0QAAAAAAMBQ6JT0OKEkAAAAupLtmnNLcSEALTst3y8Mx1VE/KeERq6tGx26LM+0fi1duRiOnRJYBAAAAAAABuA5oaTtckJZJkJJAAAAdCXjNWe2DswAdKcJteyb38FoQiG/lb2A++5s0ml5vvW7WR+UNxFxkH0SAAAAAABgCJ4TSspWOLQsJ+kBAABAVy6SzWy2DswAdKMJGMzN7WB8Ks8XrBl9WUTEcUT8u3TrYhhOdVoFAAAAAID6PSeUlK1wyGmNAAAAdC3btadQEgBtOE3Y1X+ImoO//lu6nVxnnwyqcFkCcu8sxyBMyuc9AAAAAABQMZ2SHiaUBAAAQNeydejNdm8BgPY13U72zGv1PpWOVmfZJ4IqnUTEL7omDcJ+RBxlnwQAAAAAAKjZc0JJ2R70ZisMAwAAYPOyHYgxKQXKAPAS2yVMQL3WuyMtrBMVu9Y1aTDmriEAAAAAAKBeTw0lZTzJWKckAAAAurZIeEK7bkkAvNRpCbhSpwvdkRigJuj4b12TqjYpn/8AAAAAAECFhJLud1HjoAAAABilbIdiCCUB8BLHCbv5D8lvETHTHYmBuizv398tYLX2yvcAAAAAAABQGaGk++mSBAAAwKZcJpvpWQVjAGBYtks3E+pzVbrMzK0NA7cooZf/RsTSYlap+R6YZp8EAAAAAACojVDS/bIVhAEAANAfnZIA4HGnETExR9X5WMLG7qczJmdlv3plVaszKd8HAAAAAABARZ4aStpLtmg6JQEAALAp18lOY5+UjhcA8BRHCe9PD8FvZW0W2SeCUbouwaSPlrc6+xFxkH0SAAAAAACgJk8JJWUrFLrxIBUAAIANy3Y4hlASAE8xjYi5mapKE6T+t3UhiSZ496vFrs68fD8AAAAAAAAVeEooaTfZQumSBAAAwKZdJpvxWQVjAKB+89JhjzpclWBxtn0LuZ2WIF6mzqa124qIk+yTAAAAAAAAtRBK+p4HqgAAAGxatgMyst1rAOD5mgDroXmrxseyJovsE0FKlyWQd2X5q/HGNQUAAAAAANTh5yeMItvpxUJJAAAAbFq2a1EFhAD8yNwMVeOdriTwJZA3K52T9k1HFeY6sAIAFWjuc07XhnHf/uTu/81TLR64b7x+wNV1+QEAgNewrwVe5V9///33j/7/mz/yrUTT/K8KxgAAAEA+rr95ieaG8Gcz14oxFN3/8EYfT3KhyLl3xxHxPvkc1OLXEsIAvjnVya0aPqMAgK5M14ouVwcsre4VbFd6H/eqFHyuF32e3/kNAEAu9rXARvwolNR8CP0v0VJcOa0ZAACAnmQrbvyPm4atEEpqj1ASK0JJ/ZqWoO4k8yRUYBkRB76r4UFHEfHB9PRuWYonFsnnAQB4ud2yn9hdK9bcG+l8LktR5+oU+nMn0gMAjIZ9rX0t9OrnH/yPZwvo3NceDgAAADbhMlkoaVehMwD3mAsk9W5Zgnnul8PDVt15BJP6NSmh8uPMkwAAPMnqZPjZWrHmTrKpm5TC1FVx6tu1/+5irbDz0n1bAIBq2dfa10KVhJJu8+EDAABAX7IV/m5XMAYA6jJLFtCtkUASPN0qmCRM2a83ZQ3GehLq+YhPte2CjrzU5OROYRSPG0P3YuqyKtRc/d6yPo/au2fPsSrovFw7fR5ewp72eexpqYk97fPY09IF+9rnsa+FnvwolJStQMgHDQAAAH3J9pAp20EoAPyYB7b9uoqIA/fJ4VlO1x5mCyb157QUZQAAec3WfoQf2nG3oPOm7HvPFXMCAHTGvrZ99rWwATol3eaUAQAAAPp0lai9ulASAOuOPGDr1VV5yLlIPAfwUpfl70cwqT97a2sAAOSwu1asuW/NN2KrdDdedTheFXOeld+uJwEAns++dvPsa6EDQknfXNUyEAAAANK6TBRKago2p27qAVDoktQfgSR4PcGk/jXdkrazTwIAjNxB+ZmVQkL6dbeY86IUcp45bR4A4FH2tXWxr4UW/PTIP2Ka7MHJZQVjAAAAILdsN7V0SwIgSiDJg7d+CCRBe1bBpKU57cVW6boHAIzHtHy/n5Vrlj9KoaDrxzo13SvfR8RfZW88d/8XAOAL+9phsa+FF3gslJTtD0goCQAAgL6dJ1sBN+8AaB7GHaefhX4IJEH7BJP6NS/fKwDAcK0XbP4vIj5ExL5ulIOzExFvIuLPchDXXFdLACAZ+9pxsK+FJxJK+kYoCQAAgL5luzZ1ww6AYw/herEsD0QFkqB9q2ASmzcRdAWAwTqIiNM7BZuMw1Yp5FydNH8sSA4AjJh97XjZ18IjHgslZSsMEkoCAACgb01h8E2iVdApCSC3bcXjvViWwIR74tCd5u/rV/PbC8UAADAc2+Wk8eae6B8RcWjtRq85af59KdI9K0W7AABDZ1+bj30t3KFT0lc3ToQEAACgEteJFkIoCSC3E12SNk4gCTbnVDCpF7olAUD9jso1yV/lpHHXhTntl6Ld63J/QFd9AGBo7GsJ+1r4Sijpq0wFXwAAANTtPNH6uDELkNe20wJ7cSSQBBvVBJPemfKN0y0JAOqzfnr8h3KyODS2IuJtKeY9LQdpAADUyr6Wh9jXktpjoaRMhUGZCr4AAACoW7aDM9yMA8jpxLpvXNOx5SzZa4YaNJ93H63ERk1KcQgA0L9ZuQ5xejxP0Rxe8rkcpnFkxgCAitjX8hz2taTzUCgpW0GQkyEBAACoRbZrVO3LAfLRJWnzfi8n8wH9aB48X5j7jTp0rQEAvVp1aW0K8fYtBc+0UzoPXOuCCQD0zL6W17CvJY2HQknZbtJnO4UaAACAegklATB2uiRt1sfysAvo10FEXFmDjfJ9AwCbd1RqcD6UAjx4ja2IeF/eUyeKOAGADbKvpU32tYyeUNJXOiUBAABQk0zFirsVjAGAzdElabOuBJKgGotSzLC0JBtz6AE/AGzEtBTWLUrR5pZpp2WTiHiriBMA6Jh9LV2zr2W0HgolZSoIciodAAAAtcnU0deNNoBcdK3YnGXpzLLI8oJhAC7L3yWbI5gJAN1ZFW1el8K6ibmmY4o4AYAu2Neyafa1jM5DoaRMb+5MhV4AAAAMQ6aOvnsVjAGAzdAlabMO3P+GKp1HxG+WZmOOPdQHgE4clXuYijbpw90iTgCAl7KvpU/2tYzGQ6GkTAVBmQq9AAAAGIZs16qKBAFyOLLOG/NbCT4AdZpHxEdrsxET3ZIAoFVHpWDuQ0RsmVp6tl7E6Z4DAPAc9rXUxL6WwbsvlJStEEgoCQAAgNoskq3IbgVjAKBbU0XhG/OpBB6AujWfiVfWaCN0SwKA15uVgw8UbVKjrfLePC/vVQCAh9jXUjP7WgbrvlBStkKgbIVeAAAA1C9bZ4PtCsYAQLeOy0lvdOvGKXowGIvy97q0ZJ1rvn8ORv4aAaArzX2704j4HBF7ZpnK7ZX36qlQOgBwh30tQ2Jfy+DolJSv0AsAAIBhuEm0TkJJAOMnKLMZBw7igkG51EVuY06SvE4AaNNJ2a8cmlUGpnnPXttrAwCFfS1DZV/LYGTvlJSpwAsAAIBhuU60Xtm6NgNk0wSStqx6534rD1aBYWlOu/xkzTq3JSALAE82K/cm3+p4y4A179335Tp5ZiEBICX7WsbAvpZBuC+UlOl04kwFXgAAAAxLpqJiLccBxs0Jbt27iIj52F8kjNiRg/Q2QigJAB7X3KM7i4jPDpZgRHbKe3ruPjQApGFfyxjZ11K17KEkp0YCAABQq0WildEpCWC8ZuVBCd1ZRsSB+YVBWwjMbMSeaw8AeNBxOdh33xQxUm+cLg8AKdjXMnb2tVQpeygpU4EXAAAAw3KeaL20ywcYL12SunfkXjeMQrP//91Sds73EgDctl32Ie/doyOBLafLA8Bo2deSiX0t1bkvlJSpVV2mAi8AAACG5TrZejmxHGB8tp1G2LlPEXE28tcImTSBmSsr3qlDD+oB4B/H5YTtPVNCMk6XB4Bxsa8lK/taqnE3lJSpS1I4PRIAAICKZQslKQwEGJ8ja9qppTmGUfJ33T1zDEB2TpGH26fLAwDDZF8L9rVUInso6bKCMQAAAMBDbhLNjE5JAONzbE07deTgLRil5tnVO0vbKd9PAGR24BR5uGV1urz70wAwLPa1cJt9Lb26G0rKdCrxsoIxAAAAwGMydUvSKQlgXI6cTNipTxFxNuLXB9nNkx1QsGnN6aGzXC8ZAL7cezuNiD9cq8F3dkqXBR01AaB+9rXwMPtaenM3lJQpHadLEgAAALXLdO2arXszwNh54NGdpfmF0Vv4O++c+QUgk91yn/HQqsODmqLmD6XI2QFaAFAn+1r4MftaepG5U1Km06YBAAAYpkWidRNKAhiP5jN9z3p25iTZHgGyak60/Gj1O3PooTwASRxHxJ+lUyDwY4dlL57pYG8AGAL7Wnge+1o2KnOnJKEkAAAAapepU5KCQIDx0H2iOxcRMR/riwO+c1y6o9EN31cAjNm0nIz93irDs+2UAs4DUwcAvbOvhZezr2Vj7oaSMhFKAgAAoHaZuiDsVDAGANqhyLs7x2N9YcC9FqU7Gt3wmQrAWO2WwrNDKwwvNomIP+zHAaBX9rXweva1bIROSQAAAFCvTJ2SABiH5rS1LWvZiY/2BpBS0x3tytJ3YivZs1EAcjgohZsOAIJ2vI2IM53+AWDj7GuhXfa1dOpuKGmSaLqFkgAAAKhdpk5JjVkFYwDgdQ7MXyeWOnpAav7+u6O7HwBjclxOwM5U+wObsF+KohVwAsBm2NdCN+xr6cx6KGk72TQLJQEAADAETkUHYCiahxiHVqsT84RhZeCb5kHxJ/PRCaEkAMbiNCLeW03ozE6pNdNpEwC6ZV8L3bKvpRNZQ0nLCsYAAAAAT5GpADnbgSkAY6NLUjduIuJkjC8MeBbdkrox8f0FwMA1h0NcOiACNmJSDgzQ8R8A2mdfC5tjX0vrfko6pZcVjAEAAACeIlOnX6EkgGFT1N0NgSQgynXBOzPRCd9fAAzVbikk27GCsDFNAednHTcBoFX2tbB59rW0aj2UJO0GAAAA9ckUSgJguJpTDPetX+suIuJ0ZK8JeLl5RCzNX+uEkgAYIoWb0K8PCjgBoBX2tdAv+1pakbVT0nkFYwAAAICnWCSaJQemAAyXBxbd0CUJWLcowSTaNRFMAmBgZqXuZWLhoFcf7M8B4FXsa6EO9rW82nooaWo6AQAAoDqXlgSAARBKat+FA7aAe+iW1A2hJACGorn2+qxwE6rxRodjAHgR+1qoi30tr7IeStpNNJUKugAAAKA+DkwBGKbtiNixdq3TJQm4z8LnQyeEkgAYgqNygjVQl0MFnADwLPa1UCf7Wl7sp6RTt6hgDAAAAPAUmQ7WUNAOMEwKudunSxLwmKZb0o0ZatXE9xkAlVO4CXVTwAkAT2NfC3Wzr+VF1kNJ24mmUCgJAACAoXANC0DtZlaodbqgAD8yN0OtE0oCoFYKN2EYFHACwOPsa2EY7Gt5tvVQ0lai6ct0yjQAAADDt0y0hpkOTQEYg2lE7FvJVumSBDzFabLrhE0QSgKgRgo3YVgUcALA/exrYVjsa3mWn0wXAAAAVC/T4RpCSQDDooC7fbokAU+x0C2pdRPd/wCojMJNGCYFnABwm30tDJN9LU+2CiVlKvi5qWAMAAAAAABjIJTULl2SgOeY65bUOt9rANRC4SYMW1PAeWwNAcC+FgbOvpYnyRhKuq5gDAAAAPAcma5lpxWMAYCn01GiXU6cA55Dt6T2CSUBUAOFmzAO78vfMwBkZV8L42Bfyw/9ZIoAAACgeplCSbsVjAGAp2kKtyfmqjU3QknAC/jcaNdWssMcAaiPwk0Ylw8KOAFIyr4WxsW+lkdlDCVdVjAGAAAAAICh0yWpXbqdAC/RHGDw0cy1SrckAPqy67oARmnuMC4AkrGvhXGyr+VBq1BSpofHiwrGAAAAAM+RqVMSAMOhaLs9S91OgFfw+dEuoVsA+tAUdp3rRgujNCl/3wo4AcjAvhbGy76WB2XslAQAAABDkymU5AYWwDBsR8SWtWrNqQO1gFdoHgRfmcDW7I/kdQAwHFOFmzB6k3LtP7XUAIyYfS2Mn30t98oYSnK6NAAAANTLzSuAYdBFol3zMb0YoBc+R9rlew6ATVG4CXnslL93ABgj+1rIw76W76xCSduJpkYoCQAAgKFxLQtAbQ6sSGsufNcDLWhOp1yayNb4ngNgU05LQReQw075uweAsbGvhVzsa7klYygJAAAAhkahMgC10UGiPR7aAG3xedIe33MAbELT6XDfTEM6hxFxZNkBGBH7WsjJvpZ//GQqAAAAgIrsWQyA6u1GxMQytWIpRAC0yOdJe5qTPqdjeTEAVKkp3HpjaSCtD+X+CgAMnX0t5GZfyxcZQ0nnFYwBAAAAAGCodI9ojwAB0KbLiLgyo63xfQdAV3ZL4RaQ27kgPAADZ18LhH0tsRZK8kYAAACAuikuBKAWirTbI5QEtG1uRlvj+w6ALkwdpgsUTRfqM5MBwEDZ1wIr9rX8E0raMRUAAABQtYXlAaASirTbcVO6mgC0ycPf9vi+A6AL56VgC6CxFxEnZgKAAbKvBdbZ1yb3c7KXv6xgDAAAAMDjtiPi2hwBVGnXg8bW6GYCdKE5zOBTROyb3VdzqCMAbZv7fknlYu3FXj/zfud2+VlxLT5ub0tht24TAAyFfW0u9rU8lX1tYtlCSU6dBAAAgPoJJQHUS9eI9uhmAnTlTCipNTMP0QFoyUFEvDGZo3KxVpR5WcLhlx13vJ+WQs7V71WRp+LO4Tsra9nl+wcA2mBfOz72tbTJvjapbKEkAAAAGKrL0vIaAPq0a/ZbcSWAC3TorJxY6wH+6wklAdCGpiDr1EwO1rLcmz0vvy97vJ5brO1N7h50sSrknJVr95n94KBMypo6DAaAmtnXDpt9LZtgX5vUzyVlCAAAANTNSTIA1MBDhHZ4cAt0aVEe/B6a5VfzvQdAG84U0Q3KshRInq8VbA7B6nT79UD1qphz9bOVfXEr1xxKdlwOGACAGtnXDot9LX2xr03oZydbAgAAAADwBFMPelpz9+Q/gLadCyW1wnNUAF7rJCJ2zGL1rsp12tmAijWf4rocirE6GGN10vyR92W1TgZWNAxAHva1w2BfSy3sa5P5Kdnr7avNHAAAAPB0ujoD1Elhdjuu3KsGNkD4sR2TchIrALxEUyT31sxVq7k2+y0ifinXuycJCuYuy2nlzev9v4j4NSIuKhgX30x0VwagQva1dbOvta+tkX1tMkJJAAAAQG0UvQPUaWZdWuEhDLAJi4j4ZKZb4foEgJeY2vtX6SYifl8r2JwnriValPforMzHb2V+6N9OKSYGgBrY19bJvvYb+9p62dcmki2UBAAAAEPloA0A+iaU1I7zMbwIYBB0S2qHUBIAL9EUXm2ZuWo0p6b/t3RAPHav9TvXpZC1mZ//RMTHysaX0Vv7UAAqYV9bF/vax9nX1se+NgmhJAAAABgGNxQB6JuHBq/XnM53OfQXAQyGEGQ7hHIBeK7mu+ONWavCx3Ja+kxg+8maPeRRmbfm9P3lQMY9RrpS8P/s3e1RHUm2LuC8ivMfrgVwLIBjAYwF0lgAbUEzFkhtQdMWCFkwyIIBCwYsGLDgggXnRkm5uxFiQ+1dX5m5niei48T5NbWzUNVbVWutBFiaXFsOuXZzcm055NoANCUBAAAAAPCWbqrcjlUazMdCYE7dYINbKz6YplwANrGr4GpxXbHhbyml/5uLEA172s5dnr6/n9dTEef8DvI5AIAlyLXLk2vHIdcuT64N4J0X6QAAAAAAvGHfAo3CriXA3Fx3httxHwRgA59SSnsWbBGros39fB4eAq7BFB7yeiriXMYnWRSAhci1y5FrpyHXLkuubdy73M0ahS5RAAAAAIDNHVuzUWgOAOZmh7ZxGPIIQB/dc9OvVmoRX/L9WtHmdJ4XcTKPHbtUALAAuXY5cu305NplyLWNexfs92pKAgAAAADYnGLs4a59RAQWoBlyHO6DALxlV4HVIrrnrP9JKZ2qCZrNqojzv1NKX4P85qUdpZQ+xF4CAGYk1y5Drp2fXDs/ubZh0ZqSAAAAgPIp+AMoz75zMpjGAGApPqoP5xkFgLecpZT2rNJs7lNKf89T/G+C/ObS3OWCwr/l88G0znOROABMTa6dl1y7PLl2XnJtozQlAQAAQB0iTUTyEgqgPAfOyWCakoCluP4MpzkXgNd094mPVmg2f+SG4csgv7d0V/l8/BF9ISa2l4vEAWBKcu285NqyyLXzkGsbpSkJAAAA6mCbdgCWYneIcWgKAJZiyupwmnMBeM2F1ZnFfZ5e3hWwPQT4vTV5yOflf0yXn9RHzfIATEyunYdcWy65dh5ybYM0JQEAAAAA8BofBoa7rv0HAFXTFDkOTboAvORDSunIykxuNUVerinbjenykztv/PcBsBy5dh5ybR3k2unJtY3RlAQAAAAAwGsUYQ/nAyOwNM2Rw2nSBeC5XYVUk3tMKf3dFPmqrKbL/z2fP8b1PqV0bE0BGJlcOz25tj5y7bTk2sZoSgIAAAAA4DWakoa7qf0HANXTHDmc+yEAz3UFantWZTK3+f572ejva91lPn+30RdiAp+a+0UALE2unZZcWze5djpybUM0JQEAAAAA8JpdqzOYZgBgaZojh7NTEgBP7efiTabxJRf+3Vnfqt3l8/gl+kKM7CildNrULwJgSXLttOTaNsi105BrG6IpCQAAAACA1xxZnUHuU0oPFR8/0AbNkcNpSgLgqW6i844VmcQvCtOac5rPK+MxVR6Asci105Fr2yPXjk+ubYSmJAAAAAAA1rFL0nB2JwFK8JCbJNneobUDIOvuCScWY3SPKaX/SSldNPa7+K47r3/L55nh9hQ5AzACuXYacm3b5NpxybWN0JQEAAAAAMA6CrCH05QElML1aBhTgwFYObcSo7tNKR3LK827yudZAec4TJUHYCi5dnwmRPpoAAAgAElEQVRybQxy7bjk2gZoSgIAAAAAYJ19KzPYVeXHD7RDMcRwmnUB6ArPjsKvwrgUbsZykzPVbfSFGIGp8gAMIdeOT66NRa4dj1zbAE1JAAAAAACsoylpOB8ggVJokhxut/YfAMBgJjiPa1W4+dDSj+JNd/m8K+AczjUJgG25h4xLro1Jrh2Pa1LlNCUBAAAAALCOpqRhHn2EBApy52QMZqckgNhMkx/Xl3xv9cwU04MCzlGYKg/ANuTaccm1scm145BrK6cpCQAAAACAdTQlDWOXJKAkmpKGs1MSQGwmN4/ni4IzFHCOxrUJgE25d4xHriXJtaNxbaqYpiQAAAAAANZRfD3MVc0HDzTp2mkdxE5JAHGZJj8ehZs8pYBzOFPlAdiEXDseuZan5Nrh5NqKaUoCAAAAAGCdAyszyEPFxw60yW5Jw2jWBYjLxOZx3Coy4wUKOIdzjQKgL/eMcci1vESuHc41qlKakgAAAAAAYBo31hUojKakYfZrPngAtmaa/Dhu81rCS1YFnI9WZyvdVPkPFR43APOSa8ch1/IauXYYubZSmpIAAAAAAHiJj2rDaUoCSnPljAyyV/GxA7A9k5qHWxVu2k2W1yjgHOas5oMHYBZy7XByLX3ItcPItRXSlAQAAAAAANPwYRIojesSAGzm0DT5wbpCvFM5hJ5uTEbf2pEBMwC8Qq4dTq5lE3Lt9uTaCmlKAgAAAADgJftWZZDrio8daJcd3IY7rP0HALARE5qHO5ZB2FC3u+cvFm0rpxUeMwDzkGuHk2vZlFy7Pbm2MpqSAAAAAAB4iaYkgDY9Oq+D7FZ87ABspnsmOrFmg/yicJMtXaSUvli8jZ14nwPAC+Ta4eRatiXXbkeurYymJAAAAAAAGN+VNQUKpYACAPoxTX6YL7kAD7bVTUe/tXobM1UegOfk2mHkWoaSa7cj11ZEUxIAAAAAAC8xgQygTQ/O6yDHFR87AP3tKoAa5Nb6MZIPdvrcmH97ADwl1w4j1zIWuXZz/u1VRFMSAAAAAAAv0ZQ0jJ2SgFLZKQkA3tYVjO1Yp6085vWDMdwpRtzYnn+DADwh125PrmVMcu3m5NqKaEoCAACAOigMBwAAAIB5fLLOWzvNBXcwlsuU0h9WcyMKXgFYkWu3J9cyNrl2c3JtJTQlAQAAQB0iNSU9FHAMAKS0aw0G8bESKJWdkoYxMAKgfcd5IjOb+5IL7WBsZymlW6va23u5FQC5dhC5lqnItZuRayuhKQkAAAAojSJJgDIcOA+DaEoCSmUIwDA+ggO0zyTm7dznAjuYin+bm/lQ08ECMAn3zu3ItUzNv83NyLUViNaU5CMBAAAAAAAAAAAv6XaMPbEyWznV/MzEumFWv1nk3hRTA8Qm125PrmVqcu1m5NoKvAt24dSUBAAAAADA1G6tMFCwKycHANYygXk7f8gYzORT3r2At+2llA6tE0BYcu125FrmItf2J9dW4F3utgMAAAAAAMZhiiJAu3adW4CmmcC8ucdcUAdzObXSvbmmAcTlHrA5uZa5ybX9uaYV7l30BQAAAAAA4CcmjgHAyw6sC0CzDl3nt3JmMAMz63Yv+GrRe7FLBkBMcu125FrmJtf2J9cWTlMSAAAA1GHfeQJgRnaBGMaHS6B0t84QAPzElOrNXaeULmo7aJpwlncz4HU7CjgBQpJrNyfXshS5th+5tnCakgAAAKAOmpIAoB43zhVQOM2TAPAzBU6b+1TbAdOMu5TSudPZi2sbQDyu/ZuTa1mKXNufa1vBojUlKeACAACA8inkBgAAAGBOxymlPSu+kS8ppauKjpf2nJsq34viTYBY5NrNybUsTa7tR64tmKYkAAAAoDSmtgMAAAAwp1OrvTHT5Fla9x75zFl4044CToBQ5NrNybUsTa7tR64t2DvThwEAAAAAAAAACExh02a6afJ3NR0wzbpIKd07vW9yjQOIwzV/M3ItpZBr+3GNK9Q704cBAACgCrtOEwAAMBJDC4fZr/ngAfjJhzxxmf5Mk6ck/h7fdlz6AQIwCrl2c3IEJfH3+Da5tlDvoi8AAAAAVOLQiQJgRu47wyj2B0pnaOEwmpIA2qKoaTOmyVMaU+XftuddD0AIcu1m5FpKI9e+Ta4tVLSmJH+EAAAAUD4vfwGWZ4e+YRT7AwBAPT44VxsxvZsSnTsrbzot/PgAGE6u3YxcS4nk2rfJtQWK1pRkW0IAAAAon6YkAAAAAOZwmCct049p8pSqmyr/6Oy8yu4ZAG2Tazcj11IqufZtcm2BVk1Jt9EXAgAAAApnxwoAAAAAGJcJy5sxtZtSPfj7fNNBSmm/8GMEYHty7WbkBkol175Nri3QqinpIfpCAAAAQOEOnCAAAAAAGJUJy/1dp5RuajlYQrpw2t/kmgfQLtf4/uRaSifXvs01rzDvqjracfgjBAAAAAAAAACIbd8goI0ojKN0dymlr87Sq9TNAbRJrt2MXEvp5Nq3ybWFidiUBAAAAJTr2rkBAAAAYAaKmPq7V7xJJfydvu5DyQcHwNbk2v7kWmrh7/R1cm1hVk1Jd9EXAgAAAAq27+QAAAAAwKgUb/Z3WcuBEt5lLjbmZTsppUNrA9AcubY/uZZayLWvk2sLE7EpSSEXAAAAtfEsCwAAAADjMlm5v/NaDhQUG79J4TpAe+Ta/uRaaiLXvk6uLci7ao50PAq5AAAAoFwPzg0AAAAAEzvMk5V5222wYcfU78I5fJXiTYC2yLX9ybXURq59nVxbkIhNSQAAAFCbSAM2bgo4BgAAAADapnipP9Pkqc1NLjrmZa5/AG1xXe9PrqU2cu3rXP8KsmpKugr0m3cLOAYAAADYhF1/AQAAAGA8ipf6u6zlQOEJU+XX28m7agDQBrm2P7mWGsm168m1BYm4U5I/PgAAAACA10UaZDUFH4IB2vbg/AJUT2bv56v7HpVSdPw69XMA7ZBr+5FrqZVc+zq5thARm5IAAACgNpF2Srop4BgAAKB1ClaG8dwCULfDPFGZtymAo1Z3KaV7Z28tzwMAbZBr+5NrqZVc+zq5thCrpqS7QL85UiEXAAAAbYj0LGtCFQAAAABTUrTUn110qZni4/VMlAdog1zbn1xLzeTa9eTaQkRsStor4BgAAAAAAAAAAJifoqV+boPVE9EexZvrHaSUdks9OAB6k2v7kWupnVy7nlxbiHdVHCUAAADEFumFshfCAAAAAEzJRPl+FL5Ru25HhEdncS2F7AD1k2v7kWupnVz7Orm2AE+bku4D/W5/fAAAANRkJ9DZ0pQEQAv2nUWgcKZHAhBVdw/cc/Z7UbxJC66cxbUUsgPUTa7tT66lBXLtenJtAZ42JUUq+vGhBQAAgFp4hgWA+mhKAkp34AwBEJQhtv10U7hvajhQeIPizfVcDwHq5jrej1xLK+Ta9VwPC/Cu+COchoIuAAAAahHpBcptAccAwHc+0gHAyzy3ANTNBOV+FLzRCn/L6xmoAlA3ubYfWYBW+FteT64twNOmpEgfmXXEAQAAQHkenBOAYrgmA8DL3CMB6qZepB8Fb7TC0JX17J4KUDe5th+5llbItevJtQV42pTkBToAAACUxwtlAKjPkXMGFMwzBgCRuQ/2o3iTllw7m2vZZQOgXnJtP3ItLZFr15NrF/au6KObjj88AAAAarEb6Ex5KQwAANOL9IwBAM/tWZFeTOGmJd47r7df6oEB8Ca5th+5lpbItevJtQt72pTkDxUAAADK4+UJAEu5t/KDKPoHaNOd8wpQLQNs+zF9m9YoRl7P9weAOsm1/ci1tEauXU+uXVjUnZJsWwgAAEAtIr08UdwHUBbX5WG8hwZKpXBlGPdHgHopUupHoRut8Te9nmcDgDrJtf3IALTG3/R6cu3CnjYlRXqBvlPAMQAAAEAfkXZZUNwHAAAAwFQUb/ZzVcNBwga6986PFuxFrosAdXL97keupTVy7XquiwuL2pSU/PEBAABQiQMnCgCqZCobUCrfyIZ5qPngAYKT0fsxOIgWmSr/sr0SDwqAN8m1/ci1tEiufZlcu7B3z/7nI3XP+eACAABA6SLtkpRMqwIojusyQJt8IxvGh3+AerkH9uNeR4v8Xa93WOqBAbCWXNuP+z8t8ne9nly7oOdNSZH+UN2UAQAAKJ2XJgBQL/dxoFS+kQEQlcnJb7su/QBhS3ZKWC/acDSAFsi1b5NraZVcu55cu6DnTUmR+OACAABA6SK9NLkt4BgA+NGD9RjExw+gVApXhnF/BKiToQH9KHCjVSbKr3dc6oEB8CK5th+5llbJtevJtQv6r2f/01cppaMgv11TEgAAAKWL9FJZYR9AeXzYGMbHYaBEvo8N5/4IUCdDA/pTyEWL5OD1XB8B6uK63Z9cS4vk2vVcHxf0vCkpEv8oAQAAKF2klyamVQHQmh1nFCiQ72MARKUgsZ+T/B8Qh6EqAHWRa/uRayEeuXZB7579T0ea7OUPDwAAgNJFenbVlARQHtfm4XwgBkrj+9gwtzUfPAAAvMBEeQAAWiDXLuh5U9JDoN9uSiUAAAClizTFPNI7CYBaaEoazo4kQGlcl4bx3AJQLwMDAF52YF0AqiLXArxMrl3Q86akaB+ZTYMDAACgZHuBzk6k3ZsBavLobA2i+B8ojW9jw2jYBQAAAACAJ6I3JdmmCwAAgFJFKxY0cRygTJpGhzG1EiiNpqRhNCUB1OvIuQNYy/sLgHrItQDrybULed6U1LkP8cu/84cHAABAqaIN0lD0DlAmTaPD2CkJKEn3jLHjjAyiKQkAAAAAAJ54qSkp0st0OyUBAABQqkiDNB4LOAYAXqZpdJi9mg8eaI5dkobTlARQJ8MCAF7nOglQB9drgNe5Ti4kelOSjy8AAACUKtIgDQXvAOWyU9JwduwHSuG72HCakgDqpCgJ4HWukwB1cL0GeJ3r5EKiNyX5wwMAAKBUkQoGFbwDlEvj6HCaAIBSuB4NpykJAAAAAACeeKkpKdJH5r0CjgEAAABeEmmQhoJ3gHJpHB1OEwBQCtejYe5rPniA4NwDAV7nOglQB9drgNe5Ti7kpaakaB+Zjws4BgAAAHgu0iAN08YByqVxdDgfQIBSHDgTg3huAajXrnMH8CrXSYA6uF4DvM51ciHRd0pK/vgAAAAoULQBGor7AMpmZ4hhNAEAJTCkbziNugAAAAAA8IydkkypBAAAoDzRBmgo7gMom+bR4TQDAEtzHRrO/RCgXvvOHcCrDPUGqINcC/A6uXYhLzUlda6b/+V/0ZQEAABAaaI9q0YbkAJQG82jw2kGAJbme9hw7ocA9VK8CfA6uzwD1EGuBXidXLuQdU1JkYqB3KQBAAAoTaSCwUiDUQBqZWeI4TQDAEvTHDmc+yEAAAAAADyzrikp0qQvHXEAAACUJtIADbskAZTPzhDDaQYAltQ1Ru44A4NpSgIAAAAAgGfWNSVFe6luSiUAAAAliTRAQ6E7QPlcq4fb8R4aWJDGyOHs8AoAAAAAAC/QlPRdpAnUAAAAlC1awbJp4wDl63a1e3SeBtMUACzF9Wc4DboAdTty/gDe5LkBoHxyLcDb5NoFrGtKumr6V//MhEoAAABKoSkJgBIpxh7ORxBgKa4/w3luAQAAAACAF6xrSkrBJl/6GAMAAEApou3mG20wCkCtNCUN5z00sIRu6MGOlR/MfRAAAAAAAF7wWlNSpJfr0Qq+AAAAKFekguVIA1EAaqcYe7gdjUnAAlx3xmGYAgAAAAAAvEBT0nd7KaXdEg4EAACA8CINzlDgDlAP1+xxfGjhRwBVcd0Z7r72HwAAAAAAAFN5rSnpLtiqHxZwDAAAAMS2mwdnRKHAHaAertnjsGMJMKfu+eLIig/mHggAAAAAAGvYKekvmpIAAABYWrRn02gDUQBqd+0MDnYQbFdEYFkaIcehKQkAAAAAANbQlPQXTUkAAAAsLVrRoOI+gLq4bo/jQws/AqiC6804rlr4EQAAAAAAMIXXmpIeUkqPgVZdUxIAAABLi7ZzguJ2gLq4bo/DziXAXDQljUNTEgAAEdjZGQCAFsi1C3itKSkF+8h8UMAxAAAAEFukgRmPeSAKAPXQlDSO9yml3RZ+CFC0riFpxyka7Lby4wcAgL4UbwIA0AK5dgGakn5kQiUAAABLijQwQ2E7QH1ugu2uPyW7lwBTc50Zh+cWAAAAAAB4xVtNSXfBFk9nHAAAAEuJNihDcR9AnVy/x6FZAJia68w4rlr4EQAAAAAAMBU7Jf3ITkkAAAAs5TDYykcbhALQCsXZ43ifUtpt4YcAReoaknacmlG47wEAAAAAwCs0Jf0oWgEYAAAA5Yj2TGqnDYA6Kc4ej11MgKm4vozj0TAFAAACkX0BAGiBXLuAt5qSHlJK903+8pcdlHhQAAAAhBBt915F7QB10lQ6ntNWfghQHE1J4/DMAgBAJIo3AQBogVy7gLeaklLAExOtCAwAAIDl7aaU9gKdh0gDUABa0w2yunVWR3GUUtpv4HcAZekaHneck1FoSgKGkPMAAKidTAsA9NKnKSnaC/fDAo4BAACAWKI9i9plA6BuirTHY7ckYGx2SRqP+x0whAJOAABqJ9MCAL30aUqKViikKQkAAIC5Rdu1V1MSQN0UaY9HUxIwpq5Y6L0VHcWj5xYAAAAAAHibpqSfRSsEAwAAYHnRBmQoZgeom+v4ePa8kwZGpNFxPJet/BAAAAAAAJhSn6aku2BnoPsIvFvAcQAAABBHtGLkaO8aAFrzkFK6dVZHo4kAGIvryXg04AK05dr5BACgAXItAEXq05SUAt7ITKYEAABgLvsppZ1Aq/2oKQmgCXaQGM+JQVnACD7kwXuMQ1MSAADReG8PAEAL5NoF9G1KumnqV7/tsPQDBAAAoBnRBmNEe8cA0CrF2uM6a+nHAIuwS9J4bn24Bkag6RyA2sjAwHMyLQA1kmsXoCnpZXZKAgAAYC7RBmMoYgdow1Xe/Y5xaCYAhuh2X31vBUfjmQUYw4FVBACgcjItANCLpqSXHZV4UAAAADTJTkkA1ErR9nj2NCYBA9htbVzubwDtMSUZAIAWyLUAFElT0np2SwIAAGBquwGnjGlKAmjHpXM5Kk1JwDZ2XT9G9ej+BtAkxZsAALRArgWgSH2bkjrXwU7hYQHHAAAAQNuiDcR49LIcoCl2khjXkWFZwBa6hqQdCzca9zZgDGoNAKhNtLpA4G0yLQA1kmsXsklTUrRJxj7+AgAAMLVoL/TtkgTQlq7R9NY5HZXdToBNnVmxUdklCRjDrlUszkP0BQAA2JBMWya5FoAibdKUFG0ymKYkAAAAphbt2dPUcYD2uLaP6ySltN/SDwIm1TUy7lniUWlKAmiTQTkAALRArgWgSHZKWm/HFpQAAABM7CjYAitcB2jPhXM6uk+N/R5gOq4X47o1cRgYiToDAGpz54wBz8i0ANRIrl3IJk1J3Ul6bOrXv81uSQAAAEwl4jOn6V0A7emu7ffO66jslgT0YZek8Wm0rZ9vu5Ri15kojqIkgNe5TpZDpqUUMm2ZXK8BXuc6uZBNmpJSwInGQj4AAABTifbMeW/qOECzLp3a0dn9BHiL68T43M+AsWgwL4+iJACAzci0ZZJrASjSpk1J0SYaa0oCAABgKtGeOaMNOgGIRBH3+OyWBLzGLknju1XYA4xIjgMAoHYyLQDQm52SXreTUjos+QABAACo1lGwUxdt0AlAJN1740dnfHR2QQHWcX0Y30VrPwhYlALOMl1HXwCAVxgqBjwn05ZLrgVYT65diKakt9ktCQAAgLFFfNb08gegbXZLGp/dkoCX2CVpGu5jwJhcpwEAqJ1MCwD09l9bLNVtSukg0BJ3hWLnBRwHAAAA7YjYlGSnJIC2XeQmGsb1KTcgAKzYJWl83bfPu9Z+VFCGTVKCQ2ehWFcBdy7f1m91HjYwgDxcDpmWEsi0ZZNr+5NrIR65diHbNCVdBWxKAgAAgDF9CLaa1wUcAwDT6t4b35ugObqT3PBlx0Ggc+Y6O4mLBn8TsJxda08DrjyDAEBoMi2tkGsBZvJui/+ZaJONd3R+AwAAMKLdYMM+kpe9AGFcOtWTsCsKkPJzhOvBNDQlAWMy9LRc3k/1p0YGAGKTacsm1/Yn1wLMZJumpIg3NCELAACAsUR8xow24AQgKkXd0zgKuMsi8LOzPEiPcX1NKT1Y02bsR18AiuDvsFyu9/2pkQFYjixBCfwdlk2u7U+uBZjJNk1Jdyml+2AnyAdfAAAAxhLx5aeJXQAx3AR8dzyX8xg/E1ijKwb6aHEmYZe/tuxFXwCKoICzXIbm9GeiPMByZFpKINOWTa7tT64FmMk2TUkp4E3tqIBjAAAAoA3RBl/cmtgFEIrmmWl0BSmfWvxhQC+urdN4tMsfMAG1BWUzRKGfPcXIABCaTFs+ubYfuRZgJts2JUWccGy3JAAAAIbaDzjlzi5JALHYcWI6Zz6gQkjdTqvvnfpJuGe1KeLuxJRDVivfXfQF2ICp8gDLkWlZkkxbB7m2P7kWYAaakvoT9gEAABgq4rOlpiSAWLqPoV+d80ns2C0FQrKTz3RcU4GxKXYr3030BdiAGhkAiEmmrYNc259cCzCDbZuSuhvaY7AT5MYEAADAUBF34fVSHCAeO09M57131RDKp4A7rc7l1rNKsxTQsSQ5rXwmyvcX8T0mQClkWpYk09ZBru1PrgWYwbZNSSngpOMDW1MCAAAwULQX+fdeigOEdBFwqNWcuvXdjfNzIazum9RHp38yteySpHFqc+6RLEkBcflcV/vbUyMDjMS1d3MyLUuSaevg2tqfXAswA01Jm9EFDgAAwLa6Z8qdYKsX8d0BAN9dWIfJdB9Rzxr9bcBfXEen81jRrn4PBRxDbRTQsaQjq18876o2o0YGGINMuzmZliXJtHWQazcj1wJMTFPSZmzjBwAAwLYiPlN6IQ4QVy07UNTqowIVaNqZIqBJXSqMbJqp8ixFkVs97qMvwAbUyAAsQ6ZlKTJtXeTa/uRagIkNaUq6yZPEIhG6AAAA2FbEZ0pNSQBx3aWUrp3/SdlFBdq0n1L65NxOSuNs2zT0sRQN4/W4ib4AG1AjA7AMmZalyLR1kWv7k2sBJjakKSkFLC7a0TELAADAFrrCwoNgC3efC9IBiEvR97QONC5Aky7y9yimca1oJwST5VmCIrd6uA/0p0YGYDkyLUuQaesi1/Yn1wJMTFPS5gQvAAAANmWXJAAiusxNqkznowmm0JQzE7EnV9sucwY9bMe9kSWoI6iHd1abUbwJDCXTbkemZQkybV3k2s3ItQAT0pS0OTcmAAAANhXxWfKygGMAYHm1FX/XyBpDG/btfja5e01JYSjgZG7Hdrmrionym1EjAwwl025HpmVuMm195NrNyLUAExralNTd1B6DnaA9oR8AAIANvQ+4YKZzAdA5twqTO7DO0IQLxT+T08QZh2+5zE1xW10e7Oi6kR1/4wCLkGmZm/t9feTazci1ABMa2pSUgk4+tk0lAAAAfUV8uXmbX4QDQHc/+BJ+Fab3q/fWULVuh6Qjp3BSjxo4Q9mPvgDMTg6rj2E6m1G8CTA/mZa5ybR1kms3I9cCTGSMpqSIN7XTAo4BAACAOkR8uekFOABPfbIas+gGiO0G+J3Qmq7o56OzOrnLSgcn3BRwDDXS5Mec9vPOldTF9XUzJ541gAFcc7cj0zInmbZerrGbkWsBJqIpaTsHbkwAAAD0pCkJgOjuUkrX0RdhBju56B6oR/et6cL5mkWtDbJ2oN3eYa0HTnVM2q6Td1ebM7wX2JZMuz2ZlrnItPWSazcn1wJMYIympO6D8n3AkyOIAQAA8JbDXCAcjYJoAJ6zW9I8jqw1VKXLzXtO2eS+5O+ZxHLsfDMTdQN16ibKP0ZfhA2dVXW0AG2QaZmLTFsvuXZzci3ABMZoSkpBi40EMQAAAN4ScdKSnTAAeMmVe8RsPipagSp8yo2ETO+88jW+LeAYamSqPHPYdy2vmqnym9nznAEMINNuR6ZlDjJt/eTazci1ABMYqykp4k3tfUppt4DjAAAAoFwRB1rYJQmAdS6szGwuc0EBUKbj3EDI9K7z1OCaPfg72YoCI+ZgkGndFG9uLuIAJmAcMu12ZFrmINPWT67dnFwLMDJNScMIZAAAAKxzmCctRePFNwDrdE1J91ZnFju5MclgLSjPoUb+WX0K9Fv50Z4GXWagkK1u3mFt7sS1FWBWMi1zkGnrJ9duTq4FGNlYTUkPedJYNKYRAAAAsE7EQRb3DUwhB2BaisPnc5BSOo/yY6ESu7lBc8cJm8V1I4U5iou251suU9rPeYt6de+wHp2/jZ1VdrxAGWTa7cm0TEmmbYNcux25FmBEYzUlpaBT3eyUBAAAwDoRnxl9WATgLXZLmteJRjAoyoVin1m5/qGAkykpYGuD3Qs3d2pHVoBZybRMSaZth1y7ObkWYERjNiVFLDza0ZgEAADAC6JOFtOUBEAfisTn9TF/YAWW1TUkvXcOZtPKLknJbrSD+I7LlOSrNniXtbkdBczAFmTa7cm0TEmmbYdcuzm5FmBEYzYl3QSdcCn4AwAA8FzUZ0VTuADow25J8ztPKR1G+9FQkNO8cxnzaakB9qGAY6jVjvsfEznNf1/Uz7us7ZyZKg9sSKbdnkzLVGTatsi125FrAUYyZlNSCtptqykJAACA5yJOFrv1YRGADdgtaV47+f29IhaYX/ds8Nm6z6qlXZI6dwUcQ81M/mYK/q7a8ZDfabEZU+WBTcm0w8geTMHfVVvk2u3ItQAjGbspKWK37Y7GJAAAAJ7YTykdBFyQiwKOAYB62C1pfjv5Hb7JjzCfw7xTGfNqrfFVAecwvuMytuOU0pFVbYp3Wts5y+9BAfqQaYeRaRmbTNsmuXY7ci3ACOyUNA7BHwAAgJWoz4hR3wkAsD27Jc1vL9+zNSbB9A7zv7cdaz2r1nZJWtHIu709OwUyMl1PCUUAACAASURBVBPl2+Od1nZ2PNMBG5JptyfTMjaZtk1y7XbkWoARjN2U1G0B+DXgidGUBAAAwErEF/ndx8SbAo4DgLp0kxtvnbPZHWhMgslpSFrOWaO/y2T5YRTcMZZuevaJ1WzOjUL5rZ0okgc2INMOI9MyFpm2XXLt9uRagIHGbkpKQbttdwR/AAAA8svKg4ALYfIWANtqtXi8dAfu3zCZ3dx0qSFpfl8aHpZgCMQwBkwyFtOz23UZfQEGOK/2yIG5ybTDyLSMRaZtm1y7PbkWYIApmpKi3tQEfwAAAKIOrPCCG4BtdY0x11ZvEQe5cQIYz26+rkUcVFCClgurHgo4hprtpZSOoy8Cg5ko3za5eHtHhvgCPcm0w8i0jEGmbZ9cuz25FmCAKZqSuq1WbwOelPf5YxMAAABxRRxY8agpCYCB7Ja0nBMfqmE0GpKW9Uf+Rtkqu9sNp7CIoUyUb1u3e8d99EUY4Fy9DNCDTDucTMtQMm375Nph5FqALU3RlJQCP0TYLQkAACCuwzypLhofEgEYqvtQ+sUqLkZjEgynIWlZjwEKq1puuJrLB4VFDHBoonwIhu5sb8czBdCDTDucTMsQMm0ccu325FqALU3VlBT1oqwpCQAAIK6oE+q82AZgDJ9yUTnLOMkNFQpbYHMakpbX3UMeGv+NCjiH2zFZngHOLV4Iig+Hea9mBniDTDucTMsQMm0ccu0wci3AFqZqSoq6BWB3M9ov4DgAAACYn6YkANjenQ/jizvSmAQbO8zXLw1Jy7kPdP+4LuAYancWfQHYyoeck2hf1DqXMV14ngDeINMOJ9OyDZk2Frl2OLkWYENTNSWl/PEyIh2yAAAA8XzIE+qiuQ4wkRyA+Zz7WLq4A41J0Nth/vcS8TmgJJGGQ5gsP9yeb7lsaFfjfDjO9zA7JvMDb5Bph5Np2ZRMG5NzPoxcC7ChKZuSok5KtkUqAABAPFE/ANklCYAxdY2un6zo4laNSYfB1wFec6whqQjXwYYkKuAch8nybOIsF/4Sh3ddw713rQVeIdOOw3WWTci0Mcm1w8m1ABuYuinpMeDJOPCxFgAAIJRuwthJ0FPuhTYAY7vIReYsS2MSrNcNp/uXhqQiRBsUGKkBa0pHubEQ3tLloI9WKZw7zyOj+ORZAlhDph2HTEtfMm1ccu045FqAnqZsSkp2SwIAACCAqLsk3ZpqCMBETB8sw04uFoqadeAlXSHCZytThN8CPo/cFHAMrbAzI31cWKWwnPvhdvI67tb+Q4DRybTjkWnpQ66JzfkfTq4F6ElT0jQ0JQEAAMQRtXDai2wAptIVqPxhdYvQfXT9p0Yx+ObCdOFi3KeUzgP+7of82xnOZHne8invHElM3T3/0bkf7MD7Q+AFMu14ZFreItMi145DrgXoYY6mpIg3tR3TIwEAAELYD/xCP+ogEgDm8ckH06L87sMrge3mZskTfwTFOMvFjBGZLD+eiI1t9HOoCRXZdzTv7eRBhT7YDWFyMu14ZFrWkWlZkWvHIddSI7mWWU3dlNS5CnpK7ZYEAADQvqi7BtymlO4KOA4A2vXgHWtxTnLhkI9YRHKY/+5NFi7H1+ADEhRwjudA1uAFu4r2yBR5j+ej6y0VOcz3AdeAacm045FpeYlMy1PuaeORa6mJXMvs5mhKivph4L2PswAAAM2Luktu1AEkAMyre7d8bc2LcpAbkw+jLwQhnObcu+d0F+Mx8GCIFc9i4zr3PZdnzjWikt15FhnVZ88QVOAwZ62dPJRDAed0ZNpxybQ8J9PylFw7LrmWGsi1LEJT0rR0xQIAALTrQ+ACRRPWAJjLaS5Cpxzdh6x/awygYauJwp/z3zvl+GTHVlPlR7aT/64g5dx5YiV4QuHWuK4UcFKw4yeFmyu/qvuajEw7LpmWp2RaXiLXjkuupWRyLYuZoynpIaX0Negp9lEWAACgXVF3Sbr30RCAGd0prCjW73komWm8tGQ1RVIBT3muFdF80313vS3gOFryay7YILbD3IwKT13m92CMY0cBJ4XqCjT/tWYgwWc5YRIy7fhkWpJMyyvk2nHJtZRKrmVRczQlpcC7Je258QAAADRpN3ChYuQdkQFYxrlilWK9z83K3oPTgtNcUHDgbBbJIMC/XJVyIA250GQb2r5/V7xCQ+y4dlxzKcxpjwL+S8+8k3DvHZ/ra2wyLW+Ra8cl11IauZbFzdmU9Bj0dPtIAgAA0J7I21t7aQ3AEiLfe0vXDef6tx2tqNhu/o71ec0USZb3m91af2AtxrfnPhbW6h7g+s86F4FrXaZykIumFXCytD6FmynfI+wSPD6ZdnwybVwyLX3IteOTaymFXEsR5mpKegg8SfmDf8AAAADNiTqAotul4q6A4wAgnptclE65PubztO8cUZHj/Hf73kkr1q3Cup+Yfj2NX/N3XeLYtUMePTzkAk7GpYCTpV30LNxc2ZPBRmc9pyHTxiPT0pdcOw25lqXJtRRjrqakFLgpaUfYBwAAaMpxflkTkZfVACzpUy5Op1wHucEjagM39djNO4D+K3C2r4Wd8n7WDYq4L+2gGnGhuTaUc8Wb9GTX8Gmsnh0OW/xxFGs33+9PtjjAA+/HRyXTTkemjUWmZRNy7TTkWpYg11KcuZuSom7/5wMsAABAOyIXxUUdOAJAORSnl68b1PV7nranCIYSrXZH+tXZKd5v+VzxM89m09jJa2vCcfu2Ldwhpq5w/otzP4nVlG4FnMxhtZvIkOv/iV08RyXTTkOmjUOmZVNy7XTkWuYk11KkOZuSUuCHiQM3GwAAgCbsBn7Bf5tfVgPAkrri9H84A1U4yufLhy1KYXekuly7frzqquBjq92B6dHNU7zJNtyTprOT72vHrf5AinCYn0/H2E3ko4Epo5FppyPTtk+mZVty7XTkWuYg11IsTUnzsVsSAABA/SK/lLGFNwClOM/F6pRvJ3/YuvExloV9yA32dkeqw6MP4m9SwDkt02LbpXiTbZkqP62d3Dju/s8UTnN2GnMwwWfDqUch005Lpm2XTMsQcu205FqmJNdStCWakh6D/kmc2BYVAACgepEHTkQeNAJAeU4Dv2uu0UH+GHvhPTkz288fav+ZiwKow5ldWt/0oEF3cqbFtmVX8SYjUNg9vc929mBk5/nvaopngSsFnIPJtNOTadsi0zIWuXZ6ci1jk2sp3txNSSn4ZGUhHwAAoF4fRp46U5OvigIBKMyd961VOsnnLnKjN/PYzR9q/5NSOrLmVflql9beDI6Y3md5owm7ucBG8SZDmSo/j1/zPc4wA4bYzzv2TrlT6o7BG6OQaacn07ZBpmVMcu085FrGINdSDU1J8/KhFQAAoF6RP9r4MAhAiS59PK1S94Hr9/zx+zj6YjCJ0/z3NeWHWqZxr1huI1cVHWvNFHHWbbVj3kH0hWA0psrP430uvDOtm218yH8/c1z7D7w7H0ymnYdMWzeZlinItfOQaxlCrqUqSzQl3eSPChHt+cgKAABQpf380jCiRy+gAChYNwjq1gmqUve+/F+5qMJHWcbwITcjfc7Nb9SnO4cPzltvkb+5zk0RZ50OZyzeIQ5T5eezl58VXH/pa7Vb6j9nfh44stPnIDLtfGTaOsm0TEWunY9cy6bkWqq0RFNSyv9YorJbEgAAQH0iP8tdKgwEoGAP+WPeo5NUre5D17/zx6796IvBVo7zh/1/5o/81OkfudCKzRggMR9FnHU5zflCkypT+OT5YzY7+fp7mQvzYJ3jnCWX2i31RD3YIDLtfGTausi0TE2unY9cS19yLdVaqikp8sPEex9WAQAAqhP5I40PggCU7sZHkiZ0H7v+ozmJDayakf6Vm9uo19fgAw2H8Lw2r8+5aIty7eYs8dk5YkJ37luze5+f+46D/W7etpoi/68CBhT8rtljazLtvGTa8sm0zEWunZ9cyzpyLdVbqimpu5ldB/7z8YEcAACgHqeBp5Dd+yAIQCW6D/VfnKwmaE7iLZqR2nLvI/cgV6Yaz+5jvkeZbFyew/xv4iT6QjCLc9ff2e3l/HfuGky29BT5l5zn+xGbkWnnJ9OWS6ZlbnLt/ORanpNracJSTUkpB9uoTt1MAAAAqhF5sISGJABq0t2zb52xZjxtTvLxi6QZqUld0cuHlNJD9IUYyHPb/E7y9UjzbDm6af//TikdRF8IZvNgl4nF/Gq6fHirHURKmCL/3I6MsDWZdn4ybXlkWpYg1y5HrkWupSlLNiVdBu6w3ckfWQAAACjbcfCX/7bsB6AmD/m9q8mObTnJBRlXPtCG1Q16u9OM1KSzXHzBMJEHQS7pIP/9+ua7rMN8Hj5GXgQWc553/GN+q+nydvmI5yw/G5S8g8hOronzt7kZmXYZMm0ZZFqWJtcuR66NS66lOUs2JT0En3KguxgAAKB8kXdJus0vwgCgJne5gYH2HOUPtKtz7ENY2/bzd5TuW9LnAidFMtwXhYejuVI8tJiuOOOfuYDLfWleuybJUwjPHss6yc8Hkd/hRnGcz/Xv+f5bugNZd2My7XJk2uXItJRErl2WXBuHXEuzlmxKSsH/UPdMdQQAAChaVwj5PvApsksSALXqhmH95uw1ay83qdzlbwyH0RekMR/yv+H/5AnBNXyYZXO3il1GF3kQZAl+zZPNffudxweT5ClIV0T/1QlZ1E4u6HMdbtNx/nf2rwoHFbxXwLkxmXZZMu28ZFpKI9cuT65tm1xL85ZuSoo+5cBuSQAAAOWK/szmAyAANfuUd+GgXTt5guS/84dauyfVa7Ur0l2ezhx5MEAEjworJmGoxPL2cmHJhfvRZFYFPP+0gx6FOcv3N5Z1kK/DVwYXNGE/31P/lXfNrdWJZvyNyLTLk2mnJ9NSMrm2DHJtW+Rawli6KSkF7547yhccAAAAyrKbp5RF1RVxP/ibBKByZ3k3Dtp3kHdP+n/5m0PkHFeL3fwR8+rJrkiKcdq3akjyrDG+O/e8Ypzk83EWfSFG1EoBD+26U0hflKM8uOBCPU6VVtf8/+R7ags+e0btTaYth0w7PpmWGsi1ZZFr6ybXEo6mpOVFn7wNAABQorM8fT+q6M/qALThIX8gMd0xlpM8bfZBg1JxVo1Il7mB7LNCnHDO8s5mTEPhUDm69wm/54IuU2S3d9hgAQ/t6uo+7p3fopzk68eFCfNVOH4ysKDFa76/w/5k2nLItOOQaamNXFseubYuci1hldCU1AXXrwUcx1JOdLECAAAUJ/IHlvv8ogwAWnCXPwJpTIpnZ02D0m70hZnZ/guNSO9DrQArvxl+MLlL97vi7OXrnkLOzXzI7yX+rXCTyvh3XqaTfD25ys+GlGW1e2rrO4fs5N/pefRtMm15ZNrtyLTUzL/1Msm1ZZNrCa+EpqTkI4SbOAAAQEFO80eWqKI/owPQnpu8OwdxPW1Q+n+5yOnMRL/JHOapqjd5IqRGJL7kvwmm9ZCvb5TnaSHnmcKNF+3mtbnL92s76VGjrjDrD2euWEe5QHBVVO9avJz9nA3vgu2eqoCzH5m2XDLt22RaWiHXlk2uLYdcC0/8n//93/8tZT0e8h9qRI/54vQQ9PcDAACU5C54U9J/5zWgDsf5xTPD/dZAsWwxL/oqd23KXLO6ooDfoy8CP1ntErn6Tw7a3GG+bq7+i/qth5fdagCc1WGemkvZHnOx7Xlu4IzsQy6i0rxKC8/kKRdl3QR/t1gL1+L5ueZ/98Xw6jfJtHVwHf2L6xsrrWTaJNdWxfV4fq7738m1/KCUnZJS8EnMO/5hAgAAFOE4+MvVrwpxAWjYef5IAk/t5V2UPuddfe7y9wo7Ka13nAssLvOwtX/nhr/3GpJ45laj7+xucoM1ZVvt4PfvJ5Pm9wOdsw/5XvuQJ8hHL+KhLQ92aa1G9GvxXA5d839ykt9PsJ5MW4fo11GZltbJtfWIfj2ei1z7M7mWH5S0U9J+/uAX1b0bAQAAwOKuAm2r/ZK/5+JS6mGnpPHYKYkVOyW179IHIzZ0nYuibvKH3asgC7ibP7Y+/e+ggOOiDo/5u9eD8zW709xoSX1u8z3morHpxk931JPBWKelqfIpF2b9WsBxsLnbfB2+NLxpa8e5WP+D3RVe9UvwAd5vkWnrJdMSWWuZNsm1VZNrh5Nr+5Fr+aakpqSk+Ms/TAAAgAVFb+4wLKNO0f9ux6QpiRVNSe3bze+iNVcwxG1utrjKH3XvcrFNjQ0Y+/m/w/zv4zj//z60sq3H/HfUUgFabe78G67eY77HrP6r6d/T8bOiTbvo0UdrBZy7+d+ta3HdWi2sH9tuLtRcFW267vf3t0BDL7Yh09ZPpiWaFpuS5No2yLX9yLXbk2sprikp+pQDBWAAAADLib5rQosvyiPQlDQeTUmsaEqKQWMSU1o1LK2alB6efOy9m3ky5arRKD25tu0/+U9BAWPTkFSGs5TS79EXoUHXT3btuymgGXZ1Pzl+0twqW7GtFt9LeWfTlpoL68e2+6RI/9i1fxDZ+XUybZtkWlrW6rdWubYtcu1f5NrxyLUU15SUcsiM3F1otyQAAID5dR8a/hN83f/b1u1V8iFgPJqSWNGUFIcpj5Tgdk3xzVtFOftrhpxpNGJpvnOVYTc/35noGsN1/pWribRP7yEPWxSEPG1oTS80te4q1GECrRZwnqeUfi3gOBjf45MizquKd03t4/DJf4o1x3ef17fVv58hZNpYZFpa0PIASLm2XXItY5FrgyuxKam7KX8s4DiWougBAABgfl3R3Engdf+atyCnPpqSxqMpiRXv52I5zB/aFLgADKchqSzRv7kCdWm5gPNGsVsY9092/Xi6C0gtdp8Uaa52CzmKflJncpvXm5/JtEBNWs60Sa4NRa5lW3JtYCU2JZlOndLfnnT9AwAAMC3PoZ5Da6YpaTyakljRlBSPxiSA4TQklcdkeaAmLRdw7ucCPtfjuO6fFHI+PPm/2+z8McTukwLBwyf//64izSJ8SSmdRl+EF8i0QE1ab0qSa5Fr6UOuDeq/CvzZd3lC8/sCjmUpnxQ+AAAAzKbll8N93GtIAiC4m/w+VmMSwHY0JJWpKwg5N1keYHFdDcxZSumzUxHWXv7vtQLJxxcKObd5Z7v7bDL5rh0NqnGSrxfRv1c8J9MClEOuRa6lD7k2qBKbklJ+mIjclHT05CM4AAAA09nPL0UiO/f3BQAakwC2pCGpbOe5YMi9DWBZF/l5I/p7SNbbeaG405T3eD7mAk75+kcyLUA55FreIteS5NqY3hX6q6/ypObIdAgCAABML/qz16MXQQDwp1Vj0qMlAejli+eJ4j0YRAFQjNOU0q3TAbzh87NdAZBpAUoj1wJ9yLXBlNqUlDxM/LlbEgAAANOwS1JKl/mDHgDwncYkgH6+5CIUynfuvgZQjA+uyUAPV/n7BX+RaQHKItcCfci1gZTclHThphV+YjcAAMCUPHNZAwB4icYkgNf9oSGpKt0girPoiwBQiLtcwAnwmp08UGzXKv1JpgUoi1wL9CHXBlJyU9JD/kOMzG5JAAAA07BLUkrX+YUxAPAzjUkAL/tFMWCVumGQ99EXAaAQ3aTofzgZwBsO1M39RKYFKItcC/Qh1wZRclNSMrH5G2sAAAAwPs9aKZ0XcAwAUDKNSQA/+iUXAlInu1sBlKN7L/fF+QDecCR//0SmBSiLXAv0IdcGUHpT0l2e3ByZ3ZIAAADGZZek79METaMBgLdpTAL4TkNS/boJxl+jLwJAQbrC+lsnBHjDiZ1KfyDTApRHrgX6kGsbV3pTUjK9+htrAAAAMB7PWHZJAoBNrBqTfFgFotKQ1I4zjbYARfGcAfTxux2CfiDTApRHrgX6kGsbVkNT0lWe4ByZ3ZIAAADGYZek7x/rFBQCwGY0JgERdc8Of/f80JQ7QyoAivKQC7IU1wNv6TLcoVX6RqYFKI9cC/Ql1zaqhqakZIr1N9YAAABgOM9WKV3mF8MAwGYeNCYBgTzma96lk96cT+5lAEVZDUBQwAm8ZicP9t61St/ItADlkWuBPuTaRtXSlHTpRmW3JAAAgIHskvSdxiwA2N6qMemLNQQatmpIunGSm3UWfQEACnOTJ8sDvEYB549kWoDyyLVAH3Jtg2ppSnqw7eo31gAAAGB7mnFS+ppSuivgOACgZg/5w6rGJKBFt3mgg4aktnUf/f+IvggAhemG9f7ipABvOFDs/SeZFqBMci3Qh1zbmFqakjoXBRzD0vwDBAAA2I5dkr4z7AIAxnPq4yrQmOu8Q9KDExvCp9yEBkA5LjxjAG+49p7/BzItQJnkWuAtcm1jampKujN58huTvQEAADZn0MX3lzpXBRwHALSkyxh/Tyk9OqtA5b5oSArnwTBEgCIp4ATW6ZpvPlidH8i0AOWSa4F15NoG1dSUlDTkfLPnYQoAAGAjXWHdkSXTmAUAE7nMeUNjElCrf/j2FNZNSum36IsAUKALQ3uBZx5zZjdE4GcyLUC55FrgObm2UbU1Jd3lyc7Rdc1Zu9EXAQAAoCcDLlK615QEAJPqCmD283Q3gFo85om1585YaJ98fwUo0qkCTiB7zMNQbizIWjItQLnkWmBFrm1YbU1JSTHZN91uSWcFHAcAAEDpPtgl6RvP0gAwvW6q26EPrEAl7vMHYMMLSPnZ2Y5/AOVRwAmkXCOmcPNtMi1AueRaIMm1bauxKenKZINvzuyWBAAA8CYTv79/hLss4DgAIIruA+s/nG2gYLe5idIHYFYechEnAOXpni/+cF4grF8MEuhNpgUom1wLscm1jauxKSn5o/xmx25JAAAArzrNO81Gd54/xgEA8+nuv38zoRco0JfckOQZgee6wZC/WRWAIp3lAi4gFoWbm5NpAcom10JMcm0ANTcl3RdwHEv7mFLaj70EAAAAL+p2lv1kab4VQtstCgCWcZUL/2+tP1CAx/zx99TJ4BXdc/RXCwSjkwcZw4UCTgjlN4WbW5NpYRoyLWORayEWuTaIWpuSkuKyP1kHAACAn53ZJembCxPQAWBRd7kx6Q+nAVhQN+jv2MdfejpVbAaj6ppCP1hSRqKAE2L4oh5sMJkWxiXTMja5FmKQawOpuSnJbknfneQPSQAAAHy3m5uSsEsSAJSiyyZ/zx/wAeb0NTdH3lh1enrIxWbuWTDcY/6Wf2ctGVFXK/M312lo1he7m45CpoXxyLRMRa6Ftsm1wdTclJQUV/1JFyEAAMBfumfFHevx7SWPDwQAm3PtZCqXuTHApF5gLv/IhXh2T2VTd4YiwijONIUykat8nVbACW1RuDkumRbGIdMyJbkW2iTXBlR7U9KFm9E3R7bHBAAA+OYw7yiLARYQkUaHcWhKYkp3Oa/8YZWBCd2nlP7HcD8G6orOfrGIsLVfcj0DTKW7Tu97FwDN+E3h5iRkWhhGpmUOci20Ra4NqvampAcfVP5kHQAAADwbrdglCWKyCwLUo5sw+ndDt4AJfM3Nj6YYM4YLRZywlT8UbzKThzxZ/qsFh6r9YsjYpGRa2I5My5zkWmiDXBtY7U1JKRec+XCb0p5/yAAAQHAf8k6yeD6EqDQljUNTJ3O5zBMgr604MILH/NH3g0zAyC7yhFOgny+5AR3m8pDv/3ZjhTrZhWQeMi1sRqZlCXIt1E2uDa6FpiS7Jf2lC4K7pRwMAADAzDwbfmeXJIjLjgjjcA1lTqsJkP8wfAsY4DbvjuSjL1P5lJ81gdd1/05OrRELOctFYJ4roA6PCjdnJ9NCPzItS5NroS5yLd+00JSU7Jb0px1FeAAAQFCf8g6yeC6EyDTTjENzF0s4zw0Ft1Yf2NBv+fohBzC1U0Wc8CrFm5TgIg89uHc2oGiP+d+qws35ybTwOpmWUsi1UAe5lj+10pRkt6S/nOSPTwAAAFHs5olJpHStmB5Cu4q+ACO4z+8aYQl3+d3ub1Yf6KFrYvyfPKAB5qKIE16meJOS3OTnimtnBYp0mws3vcdfjkwLL5NpKY1cC2WTa/lBK01JyW5JP9CgBQAARHKed45FQSJEd+f92GAauyjBp9xoYNckYJ3V7kg++LIERZzwI8WblOghF4cZeABluVa4WQyZFn4k01IquRbKJNfyk5aakuyW9JcjIREAAP4/e3d71Ub27Au4POt+RzcCNBGgiQAmAjMRgCMwjsAQgXEEhggGIjBEMFIEAxFcKQLu6r9LY2He9NKSuns/z1pannPOh9OqDWi3un67KMRBTozlxxc/mumBq+IrsBp/R2mK4czUJGFDYMp0JJpCEyf8oHmTpqv2DH+6p4BGuMznGSZ0N4c9LfxgT0sb2NdCc9jX8qwuhZLCtKRHqlr0GnQ9AAAA66AZ7ye1AEKoZmVCXTTNaYaTbq0MFM90JJqmalr7YFUo2FfNm7RE9T1B3z0FbNUHnxmNZU9L6expaRP7Wtg++1pe1LVQkmlJP+1ExElTLgYAAGANjnNSLKYkAT9dObRnaddO9aKh7vLUuQ9+v6FI1V7/d4cQ0FAXmjgp1AfP4mmZcd5TfLJwsFH3Oen0QtkbzZ6WUtnT0kb2tbAd9rW8qWuhpDAt6ZHPmQwGAADomp5DKR7RoAhMjU37WZq60XQX+X3vpZWCIkyyQeggw4nQVNXn05+ez1KI6d9mTTi01Xk2ko2sIKzdtUmnrWJPS0nsaekC+1rYHPta5tLFUJJpSY/ZPAIAAF10mhNi+dGYbEoSMMv3QYubqBstMc5pkX964Aqd9jVDiD6baIubDNBp4qTLJvlz7m8zbTfMhrIzKwlrU01vODSRu3XsaSmBPS1dYl8L62dfy9y6GEoK05Ie2c8/CAAAAF1Rfbn40Wr+x5Qk4FfVA/RbVVmIQ45om5vcE33yXTh0ym2e8nriQS8tNMwwndAsXTRyKjAddOp0eajdff5e+Z6pvexp6TJ7WrrKvhbqZ1/LwroaSjIt6bEq2d5r0gUBAACswP3eT9WUpLumXAzQKAKL85v4bKHFzrNZ5tIiWZBPzgAAIABJREFUQqtVD3k/5GnFmoNos3E2uflcoksu8++z71/oIqfLQ30uNft3hj0tXWRPS9fZ10J97GtZSldDSWFa0iM7GlEAAICOOMmJsPzgXg94iWlJ8zs3jYKWq35+j/PUOr/30C6TbJYY5AFz0BXHOc0P2u5T/jy7X6DrTt1PwNKqPf1fPi86yZ6WrrCnpST2tbA8+1pW0uVQkmlJj33Mh1oAAABt1RPCecSUJOAtJyr0pnufLXTIME88/TN/toFmm544eeohLx11no1APpNoo0nuqfQbUJLp/cQnBwDD3K5zevGVknWWPS1tZk9LqexrYXH2taysy6GkyA2Vm4KfnLIHAAC02UVOguUHTfTAW6oHL19V6VXHDb42WNZNPjz64PtxaKTqpNbf8zPIIQN03TDDd9dWmha5zb3UjUWjUOf5O3DpBwBedJ+nyB86YKAI9rS0kT0t2NfCPOxrqU3XQ0ljTVqP7DkhFwAAaKnqNKP3Fu8/XzUwAnM6FUp40VcPZem4i2yaOXMiJDTCbZ5QfGAvT2HG2djwycLTAp/y77RGHEo3zgD1n7mHAX76mvfaTpEviz0tbWJPCz/Z18LL7GupVddDSZEPXjVe/HSa6V8AAIC26Jn8+sjEARzAAqYPzHls5G8phRjPfCcsnATbMZoJIwnDUrLqhOI/8ncCmmaUP5/nVgYeuck9jCms8KOR+Y88DFqjf7nsaWkye1p4mX0t/GRfy1qUEEoKDQaP7Nh4AgAALVN9GbJr0f5z7sshYEHDfNDCD5M8Gc/fUkoinASbd5+fvwNhJPjPcGaKHzTF9GTgoRWBF5nCSskmua8/8FlBsqeliexpYT72tZTMvpa1KiWUdOGEgkfeOyEXAABoiepLwc8W6z8TB00AS7rIB5P8+F7Ml+2USjgJ1m+UD3f7Jr7Ci06dME8DTCfZnVgMmMvsvcSlklGIM/t6XmFPSxPY08Li7GspkX0ta1dKKClsvJ6o/rD0GnZNAAAAv/KlyGOnJnsAKzjxgOV/TeKmVYBwEqzDbTYCDdzHwFycMM82nZlkB0sb5/Th333HQIdd5s+47+N5iz0t22RPC6uxr6UE9rVsTEmhpJt8IMQPO/lHBgAAoKmq5vk9q/Ofe1OSgBocF/xw5YMmcXhiNpz0KfcbwGKmYaQDjUCwlNNsjvAcl024nWnGAVZzp4mTDpru7Y/zZxzmZU/LJtnTQr3sa+ki+1o2rqRQUpiW9MTHfEgGAADQNH1fpj+hHkBdqi+gvxZUzWoCzF8CSfCqcYaf+xngGykXvGl6yqQwEqzuLn+X/hKQZU3u8+frQDMO1E4TJ13goAHqYE/LutnTwnrZ19IF9rVsTWmhpKEPiyeqZoxew64JAADgIie88sOtZnqgZicZPOi6+/zi/coPEMyt2nMM8sHVtbLBI1XQ9Swi/q9TJmEtrjIge5a/b7Cq6d/tgXsCWDtNnLSRpk3WwZ6WutnTwmbZ19JG9rVsXWmhpHCy9BO7agIAADRM1Si/b1Eecd8GrEMVPPijwyd3XueD2mEDrgXaqHpwdZgPX79qpKFwowzz9nJvPi69ILBmp9nIWdJ0T+p3mfcD/m7DZs02cWrIp6k0bbIJ9rTUwZ4Wtse+ljawr6UxSgwl3eUHBD99zM0rAADAtvUEcJ649QUSsEbD/F6oSw/HJ9k4fuhBLdTiLkPj/fzdGikrBbnMAO/A5FLYuHF+/jiZmEVd58+NiXawXXczDfmfOnwgCu1ymZ8RmjbZFHtalmVPC81hX0sT2dfSOCWGkirnUqtPeJgGAAA0QXVvsmMlHjlu0LUA3TR9OP5HBiHb7DIfDPmuC+o3zt+tQf69uPQ9Ox11nw0G/zf34ibuwXbNnkyskZPXTE8HPtS4CY0yzh6d6l79r2yyhk2a5OHVmvvZJnta5mVPC81lX8u22dfSaKWGksZO3n5iT00AAIAtq75gf28RHvnqyyRgg4Z5otafLQwnXc58CW86EqzfMH/fptOT2h5ohMnMVKR+Nhj4PIFm0cjJSy7zHsbpwNB8V/kd8O/5vadDDlin27xf7WU/lO/ZaQJ7Wl5iTwvtYl/LJtnX0grvHh4eSl6p6hdztwHX0SR/OPUPAADYgl7eo5mS9NMkGyI1Q/Ka6gHVdxWqxZkDW544yIfkhw39+3yfU1sufAEPjdDPvxnHvnenRa6zieDKvhtaZ/q5c+K7hGJdtqwZp+jGjDm4Jy/XscOqqNEk9/bnep9oCXta7Gm7xZ62bPa11Mm+ltYpPZSkceepUUQMmnZRAABA5135gu4JX1wzD99t1Mfv3Mt6+SDloAEBpfv8zLjJf4FmGmRDTVNDjZRtlIHWK6FW6ITpXvVUKLYIk2zIaePBBBo4X+eenH7+Pa+aOfeKrwaLmh42cKFytJQ9bVnsabvLnpawr2VF9rW0VumhpMgGhv0GXEeTfM0HxgAAAJtQ3X98UelH7vMLS3iLUFJ9PCya3yBf/fy3l686H67c5r93+Rrm93imWED7HM68BJTYFtP1oAzTSZ9H1rtzRjONm21VfGPGG9yTM2swc9K85nxe4rABusqetrvsabvPnpZf2dcyD/taOkEo6UfzxL8NuI6m+TMbPQAAANapn43mGlQf+8sEEOYklFQfD4sA1k9AiU0a5XOOi7znAMrRy6YfpxK32yS/GznvyN/x4hsz3uCenJdo5GTW/cxng4ZNus6ethvsactiT8tr7GuZZV9L5wgl/VD9Un9swoU0yH1+CDp9FgAAWCfTa5+6zaAJzEMoqT4eFgFsloewrINTJYFf+bxpn9uZv+VdelatMeN17smZx2DmkAMN+uWwxwd72jaypy2TPS3zsq8tk30tnSaU9EMvf8GdzPjY14g4adIFAQAAnVLdb3yxpE/84SR3FiCUVB8PiwC2p58PYKvPtffWgQVM8qCDqw42+gD108zZXCU05mjMeJ17chbVz/uH6X2Efp9uuc7PhBsNm/CEPW1z2dNiT8sy7Gu7zb6WYggl/aQZ7nl/5R9EAACAOg3yixdfqj3mcAgWJZRUHw+LAJpj+gD2wEmRvGGUPyfCSMCinEq8faWdEKwx43XuyVnVwczLZP72Gc0cNnBTejFgAfa022dPyyx7WupgX9tu9rUUSyjpsaEN+hOTTOJ6oAcAANTJ/ddT7r9YhlBSfTwsAmim3i8PYu0h+ZVgEsuY3nv5uSFmTiWenkzsAJX1KfmEYI0Zr3NPTp2m9xADzZyNNW3WnL7syWB19rSbY0/LS+xpqZt9bfPZ10ISSnpMI8/zrvNmBQAAoA7Vl7GfVfKJTxFx3rBrovl8l1EfD4sA2mE2pDTwIJYkmMQienlQxl3+3MCvBr8EYjV0Lm+2OeeqrW+iJhozXueenHWbbeas/t1V8Y2Z5N7rZuZf+3ZYP3va+tjT/mRP+zp7WjbBvnZ77GvhFUJJT1Ubx/dNu6gG0BwHAADUQYDieaP80hAW5XeqPh4WAbSXB7GEYBJz6mXDwHTq2teIOFE83tCf+YwRiH3d7UxjjuYcoMl6v9xDuI+oz/SzYPYFbJ897fzsaYE2sa9dH/taWIBQ0lP9/MPhdIDHJvlhVdrIUQAAoD7T06h9CfbUn/lgAxYllFQfoSSA7ph9ENvP/96zvkW4NfmGV/waSJr6EBEXCseCBs+8Snu+PPqlMcf3GkAXTJs5ezP3E77Pft5t9hDd5WfAnZ4iaB17WntaoLvsa+dnXws1EEp6XtWA8rmJF7ZlTu4GAABWYTLt8y4j4riJF0YrCCXVRygJoPumDTbT04F7wkqdZH/Nc14KJE394bRTatCb+azpzYQk234K/ShPh7/5pUkHoCSzf9t7M/9zl+8nJrk/Gv/yryZN6DZ7WoBus6+1r4W1EEp62Z1U6LM06AAAAMuomgK/qdwTk2yKHTfsumgPoaT6+M4DoFwlPojtOsEkZr0VSAr3ZmzItKFz+jnTmzkQclufO5OZQN60MefulxcAb5v+je/nK2b+3kfDTqYfzex5Zhsxf/0cAHiOPS1At9nXAksRSnqZpp6X/emkAAAAYAH9/OJnR9Ge+BQR5w27JtrF9xf1EUoC4DmzIaVpk81s443gUnONcq8kZFK2eQJJU35maJLZ5p9Zs41A83iuAUdTDsD2zd5f/Opgyat7qY9naH8DbIk9LUD32dcC/yOU9LqriHjf5AvcEqfFAQAAixhq1nzW6JUv6GBeQkn1EUoCYBUXEXGkgo0jZFK2RQJJU6ZsAQAAAADAAn5TrFedZACHx3byASsAAMBbzgWSXnTS0OsCAGBxxxlmoFn2MpSyyAnMdMMygaTIcKF7NQAAAAAAmJNQ0uvunJD7ovceygAAAG+oTiT/qEjPunxl7DgAAO0kmNRMgknlWTaQNPUlIg5LLyIAAAAAAMxDKOlt1aneo6Zf5JZUD2UGRb5zAADgLVUT2JUqPWvikAcAgM6qgkm3lrdxqnDK0DONIvRXDCRNXfh5AQAAAACAtwklzUez2MuunC4IAAA8o7pX2FGYZ1X3mOMGXhcAAPU4dNhZI+1mWEXQpLsGGT5bNZAUeT974RkYAAAAAAC8TihpPtVDqq9tuNAt2M2HMgAAAFOnEbGvGs+6dQ8FANB5VQD9QDCpkXbymc9x6YXooMNc2zoPx9hz/wYAAAAAAK8TSppf1VQ3acvFbth706QAAIBUNV9+VowXaX4EACiDYFJzVaGVb55rdEq1ln+vaVpv9QzsvODaAgAAAADAq4SS5jfWPPaqLxExaPD1AQAA69eLiCt1ftFZRNw19NoAAKifYFKzfckpOL3SC9FivVzDL2t+Cx89IwQAAAAAgOcJJS2maq67bdMFb9iVh3cAAFC0qzWdTN0F9zmBFwCAsggmNdtRRNx4ttFK/Vy7ow1d/LnD+QAAAAAA4CmhpMVVJ6FN2nbRG7KbJ9IBAADlqRq09q37i5yqDQBQLsGkZtvLiaYHpReiRQ4jYphrtyk7AmwAAAAAAPCUUNLi7pxu/ar3EXHS4OsDAADqVzWEfVTXF33N5jUAAMolmNRsVeDku+cbrVAdiPH3lqb07ri3AwAAAACAx4SSllM98Lht44VvyBcnCgIAQDH6Jqa+6t7BFgAAJMGk5queb1yZhtNIg5yOtO0DMfbcAwMAAAAAwE9CSctzWt7rPLQDAIDu6+XefxsnVLfFSTafAgBAzASTJqrRWO8j4s7ha41ykhOK9hpyUUeeEwIAAAAAwA9CScurTmM7a+vFb8BOPiACAAC667xBTWFNdJ2hLQAAmCWY1HzVM47vec/jALbt6eezpi8NPAzji+AaAAAAAAAIJa3qNCJG7X4La1U1J150+P0BAEDJjvN0aJ43yRoBAMBzhoJJrfBxZq3YrOoZ3L8Rsd/gul9lcAoAAAAAAIollLQ6TWavO1IjAADonEFEfLOsrzrOE/ABAOAlgkntsGtq0kZVvxN3EfG5Bde6k8EkPxcAAAAAABRLKGl11UPDs7a/iTU7z6ZFAACg/apmqxvr+KrrbEwDAIC3DPP785FKNd50atJh6YVYk37eR33PIFhb7EXERdcWAwAAAAAA5iWUVI9TDwxf5aQ4AADojpvc4/O8iWmxAAAs6C6nw3jO0HxVWObvvC/ql16MmvTycLt/I+J9S9/D+3xWCAAAAAAAxRFKqo+ms9ftOikcAABa7yJPgeZl1b3hWH0AAFjQWDCpVfYzRHPhQLal9TLIc5dTqNrus2eFAAAAAACUSCipPsOIOOvKm1mT/XxABwAAtE/VXHVk3V517TAGAABWIJjUPkcZqjkVTprbbBjpc8cm8VYTnwYNuA4AAAAAANgYoaR6nXpY+KYjJ8UBAEDrVI2R3yzbqybudQAAqIFgUvvsZLhGOOl1/Ty4rothpKmdPKjCzwAAAAAAAMUQSqqfJrS3fXNSHAAAtEbf9J+5HGcDKQAArEowqZ1mw0kXeS9FxGHeU/6bB9d1MYw0azcibppzOQAAAAAAsF5CSfUbRsRZ197UGtx4IAcAAI3Xy+axrjeNrepacAsAgJoJJrXXToZv/s1nIYcF1qCfU6OqgNbfEfG+Ade0SXsZTAMAAAAAgM4TSlqPUw8K37STTXu9hl8nAACU7CKbqXjZxMRcAADWRDCp/fYzlFOFc84jYtDh99rLe6NhBrI+59SgUh25VwQAAAAAoARCSevjQcPbnBQHAADNdV7gadbLOM5mUQAAWIdpMOladVutCud8jIh/MrRz2pGAUvUeTvI9/b+I+OZgi0e+dTyIBgAAAAAAQklrVD2A+dTZd1ef99nsCAAANMdxNszxuq85ARYAANapCiYdRsSlKnfCXk4R+icnKF3k+vZa8Ob6eb94kddevYcvgkivusm6AQAAAABAJ717eHiwsutVPWzY7/IbrMkHU5MAAKARBtlYxuvus1amJLFt1eSE71ahFmc5tQAAmqz6Hv3ICnXWKJ8rDWde29LLe56D/HeQE59Y3Cjr6P4RAAAAAIDO+T+WdO2O88HRTsff56q+NeABGwAAlG6QDXC87VhDGQAAW3Cc/y8Fk7pp75mpQ7c5legun6GMZ/5dVT9f0wBSbyaA5LlWfao1PZ/5/QUAAAAAgM4QSlq/u3zI8HfX32gNbvKkOMEkAADYvF6euq7x7G1nwlsAAGzR9DC0LxahCPv5eslowYBS38SjrTjKZ4YmcwIAAAAA0CnvHh4erOhmXEXE+xLe6IpGGUxy4jgAAGzW8JkTuXlqlKeGQ1NU99DfrUYtzjSJAtAyVTjpm0WDVvkrnxkCAAAAAEAn/GYZN6Z6OHhfyHtdxV6eON5r71sAAIDWuRBImsskIg5bcJ0AAJSh2sd/sNbQKhcOugAAAAAAoEuEkjZnnMEk3lY1Q56rEwAAbEQ1FeRIqedS1equBdcJAEA5qoDDHxmgB5pvJyclOZwPAAAAAIBOEErarGoC0FlJb3gFR4JJAACwdtXBCZ+VeS7X7lEAAGioYUQcCCZBa+xmMAkAAAAAAFpPKGnzqpO1R6W96SV9NF0KAADWpmpa/Ka8c7l3bwIAQMNNg0meP0A77Dv4AgAAAACALhBK2o5DJxbO7ZvmPwAAqN3AqcwLqe5Jxi26XgAAyiSYBO3icD4AAAAAAFpPKGk77jxkWMh5Nk0CAACr60fETUTsqOVczrJeAADQBuMMJl1bLWiFb56BAQAAAADQZkJJ21OdSn5Z6ptf0E42AXooAwAAq+nlvYhA0nxuI+K0DRcKAAAzqmDSoWcQ0Bo3eb8OAAAAAACtI5S0XScRMSq5AAvYyeZJD2UAAGA5vWx02lO/uUxMuAUAoOWq/ewniwiNtyOYBAAAAABAWwklbdc4HwpOSi7CAnY9lAEAgKVdCCQtpLpXu2vR9QIAwHPOI+KDykDjVffrA8sEAAAAAEDbCCVt3zAiTksvwgL2BJMAAGBhVSDpvbLN7WtOaoU2GFul2qglAF1V3Q/84YA0aLTLfP4FAAAAAACt8u7h4cGKNcOVJsGFXObJ5QAAwOuqBsQjNZrbyOnUtJAvd+rxp0ZQADpuYIIqNNJtRBxYGgAAAAAA2sikpOaoAjb3pRdhAUf58BQAAHjZiUDSQqqT4w9bdL0AALCIYQYfblUNGmPkPhQAAAAAgDYTSmqOsYcOCxNMAgCAl1UHH3xRn4VUNbtr0fXC1EQlajHuwHsAgLeMM5h0qVKwdff5+2gfCgAAAABAawklNUt1SuGH0ouwoKM8/R0AAPipCtd8U4+FfI2IqxZdL8waqkYt1BGAklT3DJ+sOGzNdFKvQBIAAAAAAK0mlNQ8F04oXNiXfIAKAAD8aGoSSFrMyGEHtJwJX6u7b/sbAIAlnEfEn6YuwsZNckKSUDwAAAAAAK0nlNRMJ9kUx/y+CSYBAEAM8qAD5jc9nRraTChpdWoIQKluMhzhmQRsjkASAAAAAACdIZTUTOMM2DidcDGCSQAAlGyQDYU7fgoWciiMQAfcWMSVqSEAJRtmSOLaTwGs3QeBJAAAAAAAukQoqbmGOTGJxQgmAQBQIoGk5ZwJItARfo5Xp4YAlG6cgf2z0gsBa/TBdGMAAAAAALrm3cPDg0VttvOI+Fh6ERY0yVMdnTQHAEAJBJKWc5v3DdAV1d+Bfau5tHctvW4AWIfDDE64x4D6CCQBAAAAANBJJiU1XzUtaVR6ERa0k81Yg1ZdNQAALE4gaTn32WgJXXJlNZd229LrBoB1ucoAv2cTUA+BJAAAAAAAOksoqR0OcvoP8xNMAgCg6/oCSUuZZCBp3MJrh9fcqM7SBLoA4KlhPpu4VBtYiUASAAAAAACdJpTUDuN8+MdiBJMAAOiqXjbRCyQt7iQbLKFrhjkFjMUJJQHA86pnE8cR8Ul9YGETgSQAAAAAAEoglNQew3x4wWIEkwAA6Jpe7nH3rOzCLjWE0XHnFnhh1xFx17JrBoBNq/YYfwhAw9wmedig+08AAAAAADpPKKldLrKJjsUIJgEA0BUCScsb5Snv0GWaHhdnShIAzGeY37Ffqxe8ahpIMqEXAAAAAIAivHt4eLDS7TPUhLgUD4IAAGgzgaTlVfcC/YgYt/UNwAKqYNKRgs3lPv82AACLOYmIL2oGT1T7y0PPoQAAAAAAKIlJSe10kE11LMbEJAAA2kogaTUHAkkU5NRiz+28JdcJAE1TfYb+kQEM4IdRPn8SSAIAAAAAoChCSe00zqY6FieYBABA2wgkreaDpjAKcxcR1xb9TZOcKgUALGeY37Nfqh/8b//tMAwAAAAAAIoklNRew2yuY3GCSQAAtIVA0mq+Ch1QqBML/6YTTaMAsLLqs/Q4Iv7KwC+UqLrvPLS3BAAAAACgVO8eHh4sfrtVDXZHpRdhSZM8uc6p6QAANJFA0mpuTZilcOcR8bH0IrzgPiL6jbwyAGivfj6v2LeGFOSDgzAAAAAAACidUFI33HjQtzTBJAAAmmiQ+/wdq7OUUe7znVRNyapg452/I8/6M//GAgD1q6YRflFXOs6zJQAAAAAASL8pRCccZtMdi9vJRqSB2gEA0BACSaupmsOOBZLgf78Dx8rwxFeBJABYq2pa4x+eWdBhtzkZTCAJAAAAAIDihVBSZ0wbjSalF2JJ02DSQSuvHgCALhFIWt2h5jD4z1VEXCvHf+4j4rQh1wIAXTbMe5szq0zHfDWVFwAAAAAAHnv38PCgJN1RPQj5XnoRVvQhIi5a/Q4AAGgrgaTV2c/DU71sDN5Vm/9NbRBaBIDNGuQefU/dabHpRN4riwgAAAAAAI+ZlNQtN9mEx/K+5YMlAADYJIGk1V0KJMGzxjlBrPTpyh8EkgBgK6ZTkz7Zj9BSt/kzLJAEAAAAAADPEErqnotsxmN5gkkAAGzSgUDSym7t4eFVVTPwScElEloEgO07z2DHrbWgRc7ynv3OogEAAAAAwPPePTw8KE03VU2N+6UXYUUfNC0BALBmxxmKZ3mjbBIbqyG8qcS/OZdCiwDQOIf53buDGWiqUe4hTdoEAAAAAIA3mJTUXYf50ITlfRNKAgBgjQSSVjfJex+BJJhPadOVR4VPiAKAprqKiH5EfLVCNNDXPPhCIAkAAAAAAOYglNRd42zOm5ReiBUdCSYBALAGAkmrm2Sj2F3b3whs2HEhDcC3pqgBQKONMzz8R35uw7ZVgfY/8+fSHhIAAAAAAOYklNRtd9mAI5i0GsEkAADqdCGQVIsTJ1fD0qrfnw8dLt+lQBIAtMYwP7f/ioh7y8aWnEXEICJuLAAAAAAAACxGKKn7htlsxGqOspY9dQQAYAUXubdkNZ8cHAAru8jm364dZPI1p0EBAO1yFRH9DIc4aI1NqaZ0/R4RpyoOAAAAAADLeffw8KB0ZTh2GnstRk5bBgBgCVW4/VwgqRaXAgdQq0EGlPZaXtZJ/m24asC1AACr6WVI5KM6sib3eaCfvSMAAAAAAKxIKKksTmWvxygbnYZdeDMAAKxd1VB304GG/ya4jojD0osAa9D2xt/bvE+/a8C1AAD16ecexXMN6jLJA0POHT4HAAAAAAD1EEoqj2BSPSY5MUkwCQCA1wgk1cfUUli/g/zeYLcltZ5ko/J5A64FAFgf4STqcJk/R4LsAAAAAABQI6Gk8miKrM8kT2K+6sobAgCgVoPce+8o68rus54CSbB+1fcGJ/lq8t8vTaUAUB7hJJZxm3tbh8wBAAAAAMAa/KaoxRnnycej0gtRg6o56+8MJgEAwKwDgaTaVIcBHAokwcaMs9l3kMGfpqmaSv/Me3GBJAAoy13uAX5v6D6FZpnuGw8EkgAAAAAAYH1MSipXPx/CaJKsx1k2bQEAQNUk9634KtRjooEMtq6ff9e2PTmpajw+9/cAAJjRlH0KzXKbz2turAsAAAAAAKyfUFLZBk5vr9WlqUkAAMWrmuG+lF6EGv0VEVedeTfQfsc5uez9ht5JNeX5Il+mpQEAL+nlHqUKouyqUrGuM8QujAQAAAAAABsklEQVTPqn+CrU5zYffmqWAgAoT9U0f2Tda/Mhawo0z7Tx9yBfdTX/TrKJ9CYDiXfWHgBY0EEeFrGpEDXbd5mBNHtHAAAAAADYAqEkIk86/qYStRllc5YHYAAAZehl8/y+9a7NpzzhGmiHXh56UjUB9/MVr/xdHOVhHtVrOPNyHw0A1KWfzz6OTU/qpPs8xOLcIXEAAAAAALBdQklMCSbVa5LNWMMuvSkAAJ7oZyBpT2lqc5n3JwAAAHU4zJfJtu13nWGkq9ILAQAAAAAATSGUxKyTiPiiIrWZZE0vOvJ+AAB4rJoKchMRO+pSG4EkAABgXXoZTjo26bZVplORLkzWBAAAAACA5hFK4lcXTgus3aeIOO/YewIAKN1x7vEEkupznQ2CAAAA69afCSiZfNs8k5yGdJGHgQAAAAAAAA0llMRzBJPq58R3AIDuOI2Iz9azVqOIOIiIcYfeEwAA0A79vB+pQkrvrdnWTIPf1fILAAAbP0lEQVRI0xcAAAAAANACQkm8RDCpfhotAQDarZfTkeyT62WfDAAANEVvJqBU/btrZdbqPichCSIBAAAAAEBLCSXxmmFE7KlQre7zYeawQ+8JAKAEvWyUsj+ul0ASAADQZIO8Z5m+dqzWym4zgHTjWQkAAAAAALSfUBKv0Xi5HpOIOMlpVAAANN8g98Waz+p1n7UVSAIAANpiNqQ0MElpLrd5Tz19AQAAAAAAHSKUxFsEk9bnLCJOu/rmAAA64jgivlnM2k2yic+p2AAAQJv1M5w0mAkqlXygxX3e5w2FkAAAAAAAoAxCScxDMGl9rrPR1enwAADNcx4RH61L7QSSAACALuvn62Dmv/c7+H5HEXE3E0AaetYBAAAAAADlEUpiXoJJ6zPKYJKmTACAZqj2vlcdbRrbNoEkAACgVL2cpNSfmbDUy//ebWhNbvPfm5l/7/IFAAAAAAAglMRCBvnAaUfZajfJYNJVx94XAEDbDHJP1tSGsDYTSAIAAHjdQf5fpwGmqWmQ6VeDOZ/Z3D7zvxv/cn9288L/HgAAAAAA4EVCSSxKMGm9ziLitMtvEACgwaqQ+Lm97loIJAEAAAAAAAAAAHSMUBLLEExar+tsiB13+U0CADRMFUb6aFHWQiAJAAAAAAAAAACgg4SSWJZg0nqNMpikcRMAYL16ua/dU+e1+RARFx19bwAAAAAAAAAAAMX6zdKzpGGedj5RwLXYy+bY4w6+NwCApqiC9ncCSWslkAQAAAAAAAAAANBRQkmsQjBpvaopVN8i4rzLbxIAYEtOIuIfkz/XSiAJAAAAAAAAAACgw949PDxYX1Y1yKk+GjrXZxQRh3mSPwAAy+tlUOa9Gq6VQBIAAAAAAAAAAEDHCSVRF8Gk9ZtkMOmm628UAGBNqj3rVUTsKvBaCSQBAAAAAAAAAAAU4DeLTE2GEXGQwRnWowp8fY+IU/UFAFjYcYa7BZLWSyAJAAAAAAAAAACgECYlUTcTkzbjNqcmjUt4swAAK+hFxHlEHCni2gkkAQAAAAAAAAAAFEQoiXUQTNqMSQaTbkp4swAASxhkSGZP8dZOIAkAAAAAAAAAAKAwv1lw1mAYEQcZmmF9qtDX9zz5HwCAx04i4h+BpLWr9vx/CSQBAAAAAAAAAACUx6Qk1snEpM0Z5dSku1LeMADAC3oZkHmvQGs3ycMIhh1/nwAAAAAAAAAAADzDpCTWycSkzdnLeh+W8oYBAJ4xDcgIJK2fQBIAAAAAAAAAAEDhhJJYt2FOTBqp9NpVE6n+zskAvY6/VwCAX51GxPeI2FWZtRNIAgAAAAAAAAAAIN49PDyoAptQhWRucqIP61eFwI41igIABehnKHvfYm+EQBIAAAAAAAAAAAD/Y1ISmzLO5kUTkzajCn/9kxMDAAC66jDDMQJJmyGQBAAAAAAAAAAAwH9MSmLTTEzavNucmnRX2hsHADqrl9OR3lvijbmfCYEBAAAAAAAAAACAUBJbIZi0eZMMJl2V9sYBgM45yEDSrqXdmFHWfVzI+wUAAAAAAAAAAGAOvykSW1A1Mw4i4lLxN2YnIv7OUFKvkPcMAHTPeUR8F0jaKIEkAAAAAAAAAAAAnmVSEttWnXJ/ZBU26j6nJt0U9J4BgHYb5L7RpM3NEkgCAAAAAAAAAADgRSYlsW3HJiZt3G5OGDg3NQkAaIHTiPhHIGnjLgWSAAAAAAAAAAAAeI1JSTTFSUR8sRobZ2oSANBU/Yi4EkbaisvcIwIAAAAAAAAAAMCLTEqiKaqpPR+sxsaZmgQANFEVWB8KJG2FQBIAAAAAAAAAAABzMSmJpqkaIL9Zla0wNQkA2LZqOtJFROxbia34kPUHAAAAAAAAAACAN5mURNNUTZB/RMTEymycqUkAwDZNpyMJJG2HQBIAAAAAAAAAAAALMSmJphrkxJ4dK7QVpiYBAJtiOtJ2TXLfd1VyEQAAAAAAAAAAAFicSUk01TCDSSMrtBWmJgEAm3AaEf8KJG1NFUg6EEgCAAAAAAAAAABgGSYl0XS9nNazZ6W2xtQkAKBug5yOZI+3PaPc4w1LLQAAAAAAAAAAAACrMSmJphvn6e2XVmprplOTrkxNAgBW1MvpSP8IJG3VKPfYAkkAAAAAAAAAAAAszaQk2qQ6Tf/Iim3VJCJOci0AABZxkHuIXVXbquuckDQuuAYAAAAAAAAAAADUwKQk2qRqnvxkxbZqJyK+RcRNRPQLrgMAML9ehpG+CyRtXTV99FAgCQAAAAAAAAAAgDoIJdE25xHxISf2sD37ETGMiFNrAAC8ogqV35l22Qifcj0AAAAAAAAAAACgFu8eHh5UkjYa5LSeHau3dffZ4HpTeB0AgJ/6OR1pX022rgrzn+R6AAAAAAAAAAAAQG1MSqKtqik9BxExsoJbtxsR37PRtVd4LQCgdL2cpPivQFIjTHLPLJAEAAAAAAAAAABA7UxKou16OaFnz0o2wiQbkc9LLwQAFOgw9wC7Fr8RRrkmd6UXAgAAAAAAAAAAgPUwKYm2G0fEICIurWQj7ETEl5lJVgBA9/UzJP63QFJj3OZeTCAJAAAAAAAAAACAtRFKoiuOI+KT1WyManLV94i4yGlWAED39HJC4r8RsW99G+MyA0nj0gsBAAAAAAAAAADAer17eHhQYrrkMIMwO1a1MSbZsHxeeiEAoEMO87PdZKRm+WTPBQAAAAAAAAAAwKYIJdFFg4i40iTbOKOIOImIm9ILAQAt1s8AuMlIzTLJyaFXpRcCAAAAAAAAAACAzflNremgYQaTRha3UfYi4ns2y/ZLLwYAtEwvJ/D8K5DUOPcRcSCQBAAAAAAAAAAAwKYJJdFV4wwmXVrhxnmfwbHTbHAGAJqtmnR4FxEfrVPj3Oaed1h6IQAAAAAAAAAAANi8dw8PD8pO11WNtF+sciPdZzjpovRCAEADHeRn9K7FaaQqfH9cehEAAAAAAAAAAADYHqEkSlE11V5FxI4Vb6TbDCfdlF4IAGiAfoaR9i1GY30Q6gYAAAAAAAAAAGDbhJIoySCbN/esemNd52Sru9ILAQBb0IuI84g4UvzGmmTYflh6IQAAAAAAAAAAANi+36wBBRlmE+e1RW+s9xHxbzZE90ovBgBsSC8nFt4JJDXaKKdYCSQBAAAAAAAAAADQCEJJlGYcEYcRcWblG+1jNkafCicBwFodZ8jlc0TsKHVjXebUz3HphQAAAAAAAAAAAKA53j08PFgOSlWFky404DbefYaTLkovBADU6CA/W3cVtfE+2AcBAAAAAAAAAADQREJJlG6QTZ57pReiBapw0klEXJVeCABYwUGGffcVsfEmuV7D0gsBAAAAAAAAAABAM/1mXSjcMJs9L0svRAtUkxz+joibXDMAYH79/Az9LpDUCqNcM4EkAAAAAAAAAAAAGksoCSLGEXEcEZ/UohX2s6FaOAkA3tbPqZD/CiO1xtec5jkuvRAAAAAAAAAAAAA027uHhwdLBD8NMuyyoyatcR0RJxFxV3ohAGBGFUY6jYgjRWmNSe5pLkovBAAAAAAAAAAAAO1gUhI8Nswm3lt1aY33Of3hItcOAErWm5mMJJDUHqOcACmQBAAAAAAAAAAAQGsIJcFT42wKPVObVjkSTgKgYL2cjHQnjNQ6l7n3HJZeCAAAAAAAAAAAANrl3cPDgyWDlx1myGVHjVrncqY5GwC6qgojneTLfqV9PpiOBAAAAAAAAAAAQFsJJcHbqqk7VxGxp1atJJwEQBcJI7XbfYbfTUcCAAAAAAAAAACgtYSSYH7nEfFRvVpLOAmALuhnEOlYGKm1rnP9xqUXAgAAAAAAAAAAgHYTSoLFVCfaX2gCbrXLDJiZTABAm/QzXHtk1VrtU+5DAAAAAAAAAAAAoPWEkmBx/Qwm7atdq91mc/dN6YUAoNGEkbphlNORhKIBAAAAAAAAAADojN8sJSzsLiIOIuJM6VqtCpV9z1DSQenFAKBxDjIE/a9AUutd5noKJAEAAAAAAAAAANApJiXBaqoG06uI2FHH1qsmGJxnAzgAbMtBTkYykbH9JhFxYm8BAAAAAAAAAABAVwklwep62Wz6Xi074T6bwauw2bj0YgCwMccZYNlT8k6ows6HOWETAAAAAAAAAAAAOkkoCepTNRJ/Uc/OmOTkpHPhJADWpDcTRtpV5M74mmsKAAAAAAAAAAAAnSaUBPUa5NQkUw665TKnJ5l2AEAd+jNhpB0V7YxJTke6Kb0QAAAAAAAAAAAAlEEoCerXywDLR7XtnNtcW83GACzjIMNIR6rXOde5tqYrAgAAAAAAAAAAUAyhJFifqvH4ygSETrrPcNKV5mMA5nCcr33F6pxJ7gnOSy8EAAAAAAAAAAAA5RFKgvWqpiZdRMR7de6kSa5v1Yh8V3oxAHik2gOcZBhpV2k6aRQRh/YAAAAAAAAAAAAAlEooCTbjOIMrpiZ113Wu8U3phQAo3CDDSEelF6LjznJCEgAAAAAAAAAAABRLKAk2p59TdfbVvNPuM5xUrfW49GIAFOQ4Xz7nu22U6zwsvRAAAAAAAAAAAAAglASbV01P+KLunTeJiKsMKGlcBuimfn6uH5uGWISvOR1J6BgAAAAAAAAAAIDihVASbM0gJ+nsWYIijDKcdKWRGaATDjOI9N5yFuE+1/um9EIAAAAAAAAAAADALKEk2K7qtP3P1qAYpicBtFc/gynVa9c6FsN0JAAAAAAAAAAAAHiBUBJsn6lJZTI9CaAdjnMykqlIZTEdCQAAAAAAAAAAAN4glATNYWpSmabTky40PgM0xmBmKtKOZSmO6UgAAAAAAAAAAAAwB6EkaBZTk8p2PzM96a70YgBsWC8nIp34HC6W6UgAAAAAAAAAAACwAKEkaCZTk7iemaAEwPoc5utIjYtmOhIAAAAAAAAAAAAsSCgJmsvUJCqTmXCSyQ0A9RjkRJzqtaOmRTMdCQAAAAAAAAAAAJYklATNV53af6JpmmycngaUhgoCsJB+TkSqPlN3lQ7TkQAAAAAAAAAAAGA1QknQDv0MouxbL9IofyaqkNKdogA8qzcTRDJ5kKlR/kyYjgQAAAAAAAAAAAArEEqCdjmOiHNTk/iFgBLAT9MgUvV6ry784iynIwEAAAAAAAAAAAArEkqC9ullAEWjNc+5znBS9RqrEFAIQSTecpvhbuFdAAAAAAAAAAAAqIlQErTXQYaTdq0hLxBQArpMEIl5TCLiJPdMAAAAAAAAAAAAQI2EkqDdetlo+9k68oZRNmRfmRIBtJggEou4zH2SYC4AAAAAAAAAAACsgVASdMMgIs4jYt96ModpQOkmIoYKBjRcP0NIB4JIzOk+Io7zcw4AAAAAAAAAAABYE6Ek6JbjDCftWFfmdJ/Tky4ElIAGGcxMRNqzMMxpkvugUwUDAAAAAAAAAACA9RNKgu7pZUPukbVlQZMMKF3ldImxAgIbNJ2GVP27q/As6DbD2XcKBwAAAAAAAAAAAJshlATddZDhJBMmWNbtTEhJkzdQt/5MCOnAlD+WVE38O8nPKgAAAAAAAAAAAGCDhJKg+6pG3VPN3qzofmaCksZvYFmzISShWVZ1lgFsk/0AAAAAAAAAAABgC4SSoAy9bNo9st7U5HYmpDRUVOAF/ZkQkmlI1KX6DDo2xQ8AAAAAAAAAAAC2SygJynKQU5P2rTs1mswElG40iUPRer9MQ9otvSDU6j7DSDfKCgAAAAAAAAAAANsnlARlOs7JSSZWsA73v4SUxqoMnTY7CWnPUrMGk9y3nCouAAAAAAAAAAAANIdQEpSrmmZxEhGf/QywZqOZgJKQErTfwczL5D3W7TLDSKbwAQAAAAAAAAAAQMMIJQH9nD7wvvhKsClCStAevZkA0kAIiQ26zTDSjaIDAAAAAAAAAABAMwklAVMHGU7aUxE27H4moDTMF7Ad/ZkA0oHPBLbgPsNIF4oPAAAAAAAAAAAAzSaUBPzqOMNJOyrDlkxmAko3pmTAWs0GkKp/d5WbLZnk/uPcBD0AAAAAAAAAAABoB6Ek4Dm9iDjJl3ASTTCaCSmZpgTLmZ2CVL321ZGGuMw9hzASAAAAAAAAAAAAtIhQEvCaqoH9NCKOVIkGup0JKAkqwWP9mfDRNIgkZErT3GYYyd9vAAAAAAAAAAAAaCGhJGAeVTP7uakatICgEiWaho/6Aki0xCjDSDcWDAAAAAAAAAAAANpLKAlYxEGGk/ZUjRYZZTjpLhvgq/8eW0BaqDcTQJqGkIRFaZP7nMB4YdUAAAAAAAAAAACg/YSSgGUcZ1PxrurRUpOZSUp3M/8trERTHGToyPQjumCSoeZTqwkAAAAAAAAAAADdIZQErOIkG4w1ytMVk18CSjcZWrqzwqzBNHQ0+OVfgU+6YhpGOhf6BAAAAAAAAAAAgO4RSgJW1ctw0olwEh03mgkqjWemLAks8Zr+L69B/t3cVzU67jL3BsJIAAAAAAAAAAAA0FFCSUBdpuGkzypKge4znDScCSzN/kt39WaCRr/+u2fdKdBlTlEU2AQAAAAAAAAAAICOE0oC6tbPZuQjlYX/TENL06BS5MSlEFxqtGnQKGYCR9PJR0JH/7+9u71NI4sCMHx2G4AOYCswHcBWYHcQSnAJKcEl2B04HeAOoAPoACrI6u7eka5n7Th8DfPxPNII4jhSfA5S/uTVgffESAAAAAAAAAAAADAwoiTgWsRJcJxDESxti//YX0ZLAqbzlaHRZ+/T66irPyA07C3/e78yeAAAAAAAAAAAABgWURJwbeIkuI5d7SJJPViqBwLllaauq64VlRa/+HX63onPIVyUGAkAAAAAAAAAAAAGTpQENEWcBO20+eL60rYWP11SeZ3oI+n373xuoFXESAAAAAAAAAAAAMC/RElA08RJANA9YiQAAAAAAAAAAADgnT+NA2hYuriyjIi/IuLF8AGg1VKM9HdELARJAAAAAAAAAAAAQEmUBNyKOAkA2kuMBAAAAAAAAAAAAPzSHz9//jQhoA2mEfE9Ir7ZBgDcTAqFnyJibQUAAAAAAAAAAADAr4iSgLaZ5gtKjxExsh0AaMRLjoO3xg0AAAAAAAAAAAD8DlES0FbjHCaJkwDgOg4R8SpGAgAAAAAAAAAAAE4hSgLablxcTprYFgCcLcVIT/nZGycAAAAAAAAAAABwClES0CXLfM1BnAQAx9vlEOlZjAQAAAAAAAAAAACcS5QEdNEix0lz2wOAL+3yv5vPRgUAAAAAAAAAAABciigJ6LJZRDxGxDdbBID/ecsx0spoAAAAAAAAAAAAgEsTJQF9MM1x0jIiRjYKwMC95BhpO/RBAAAAAAAAAAAAANcjSgL6ZJzDpBQoTWwWgAE5RMRTfvYWDwAAAAAAAAAAAFybKAnoq4ccJ81tGIAe2+QQ6dmSAQAAAAAAAAAAgCaJkoC+m0bE9xwpjWwbgJ54ySHSykIBAAAAAAAAAACAWxAlAUMxjohlvp40sXUAOuhQXEXaWiAAAAAAAAAAAABwS6IkYIgecqB0b/sAdMCmiJEAAAAAAAAAAAAAWkGUBAzZNF9OSoHSyCcBgBZJV5Fec4y0thgAAAAAAAAAAACgbURJAP9Z5mduHgDc0K64irS3CAAAAAAAAAAAAKCtREkA76XrSd8j4sH1JAAa9JJDpJWhAwAAAAAAAAAAAF0gSgL4nOtJAFyTq0gAAAAAAAAAAABAZ4mSAL6Wric95kDJ9SQAznGIiNccI61NEgAAAAAAAAAAAOgqURLAcR5ynHRvbgAcYZNDpFdXkQAAAAAAAAAAAIA+ECUBnGaaA6V0QWlihgB8YFdcRdoaEAAAAAAAAAAAANAnoiSA881ynJQipZF5AgzeS46RXoc+CAAAAAAAAAAAAKC/REkAl7XMcdK9uQIMyltEPOcQaW/1AAAAAAAAAAAAQN+JkgCuY5wDpfTcmTFAL+0i4imHSFsrBgAAAAAAAAAAAIZElARwfdN8PekxIibmDdBpuxwhpatIa6sEAAAAAAAAAAAAhkqUBNCsWb6e9CBQAuiMQxEirawNAAAAAAAAAAAAQJQEcEsCJYD2qkKk6gEAAAAAAAAAAACgIEoCaIeH4hnZCcBNCJEAAAAAAAAAAAAAfpMoCaB9Upi0cEEJoBFCJAAAAAAAAAAAAIATiJIA2m0WEUuBEsBFCZEAAAAAAAAAAAAAziRKAuiOKlBKV5Tu7A3gKLsiQloZHQAAAAAAAAAAAMB5REkA3TTN15PSM7dDgA9tihBpbUQAAAAAAAAAAAAAlyNKAui+cREopStKIzsFBuxHvoSUQqStDwIAAAAAAAAAAADAdYiSAPqnipPS68R+gZ7bFRFSet1bOAAAAAAAAAAAAMD1iZIA+m1aREr3dg30xCYinnOEtLZUAAAAAAAAAAAAgOaJkgCGxRUloItcQwIAAAAAAAAAAABoGVESwHBNi0ApvY58FoAW+ZEDJNeQAAAAAAAAAAAAAFpIlARAZVYESnNTARq2qV1DAgAAAAAAAAAAAKDFREkAfKa8onRnSsCFbYpLSOnZGzAAAAAAAAAAAABAd4iSAPgd4xwnLURKwIlESAAAAAAAAAAAAAA9IkoC4BRlpDSLiLkpAjUiJAAAAAAAAAAAAIAeEyUBcCmLWqg0MlkYlLccH61FSAAAAAAAAAAAAAD9J0oC4FpmRaCUXicmDb2xK+Kj6hUAAAAAAAAAAACAARElAdCUcS1Sck0JuuOtFiFt7Q4AAAAAAAAAAABg2ERJANzSrPbMbQNubpPDozJCAgAAAAAAAAAAAIB3REkAtI1QCZpTBkhVhAQAAAAAAAAAAAAAXxIlAdAF9VApPSObg6O85fBoK0ACAAAAAAAAAAAA4FyiJAC6apqfRY6U0vs724TY1a4fVSESAAAAAAAAAAAAAFyMKAmAvqkCpZlYiZ7b5dholV+3rh8BAAAAAAAAAAAA0BRREgBDUY+VxhExt306YJODo7X4CAAAAAAAAAAAAIC2ECUBMHTjWqi0yPMQLNGkFB7tc2y0rwVIAAAAAAAAAAAAANA6oiQA+Ny4uLBUfybmxhEOOTSqB0fCIwAAAAAAAAAAAAA6SZQEAKerh0pVxBQuLQ1OdemoHhtVERIAAAAAAAAAAAAA9IooCQCua5ZjpTJYKr92Z/6tVsVGySq/lteNVh37eQAAAAAAAAAAAADgIkRJANAOZbRUXV6K2tcjvx/Z2cneij+4LoKjMjQq3wMAAAAAAAAAAAAAHxAlAUC3LWp/++oKU6n+PZV5R37y8lpRaf3B1+uXiz76HgAAAAAAAAAAAADgTKIkAOAz5cWma3GVCAAAAAAAAAAAAAC6JiL+ASIGZFTrDc8HAAAAAElFTkSuQmCC"/>
</defs>
</svg>
